     M  2   �  2   ���`$f\FWG��Љ@            '      >      Q      X      c      r      y      �      �      �      �      �      �      �      �      �                1     8     [     ~     �     �     �     �     �     �     �     �          ,     ;     B     U     `          �     �     �     �     �     �     �     �     �     �               "     )     0     7     >     I     X     c     v     �     �     �     �     �     �     �                    #     *     y     �     �     �     �     �     �     �     �     �               %     4     ;     v     �     �     �     �     �     �     �     �     �     �               9     H     c     n     }     �     �     �     �     �     �     �     �     �     �     �                +     :     E     L     _     n     y     �     �     �     �     �                    $     +     6     A     H     S     ^     e     x     �     �     �     �     �     �     �     �     �     �     �     	     	     *	     E	     X	     _	     j	     �	     �	     �	     �	     �	     �	     �	     
     
     
     
     *
     E
     P
     _
     j
     q
     �
     �
     �
     �
     �
     �
                    #     .     5     @     G     R     ]     l          �     �     �     �     �     �     �     �     �               /     :     E     T     _     v     �     �     �     �     �     �     �     �     �     �     �               0     7     B     a     l     s     ~     �     �     �     �     �     �     �     �     !     0     ;     J     ]     d     o     ~     �     �     �     �     �     �     �     
          $     ?     R     e     l     s     �     �     �     �     �     �     �     �     �     �     �     �     �     	               .     =     H     S     j     u     �     �     �     �     �     �     �     �                     !     0     ;     B     ]     d     s     z     �     �     �     �     �     �     �     �     �     �     �     
          $     /     F     Q     h     s     ~     �     �     �     �     �     �     �     �                          +                     �                  �   +              ����   �      *            �   �            	      �   �         
      �����   +  
            �����   �                �����   �   	               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                      �����   �      	         �����   �                  ����                        ����                        ����                        ����                            +      "               �               �����   +           	         �         
      �����   �                  ����                        ����                     ����   v               ����w   �                  ����                        ����                        ����                        ����                        ����                        ����                            +                     �      !         �����   +     +      	         �         
         �   �                  ����                        ����                     ����   �                �����   �                  �   �      *         �����   �                  ����                        ����                        ����                        ����            2         �����   �               �����   �                  ����                        ����                        ����                        ����                        ����                        ����                            +                     �                  �   +      $      	         �      2   
      �����   �               �����   �   !            �����   +  "            ����   �      2         �����   �                  ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   #            �����   +  $               ����                        ����                        ����                        ����            #                +                     �   %   #         �����   +  (   #      	   ����   �   &      
      �����   �   '               ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   )               �   +  *               ����                        ����                  	      �   �   +      
      �����   +  .   *         �����   �   ,             �����   �   -               ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   /   "         �����   +  0               ����                        ����                        ����                        ����            "                +      +               �   1               �   +  4   +      	   ����   �   2   +   
      �����   �   3             �����   �   5   "            �   +  6               ����                        ����                        ����                        ����                        ����                        ����            "            �   �   7               �   +  :             �����   �   8             �����   �   9   	            �   �   ;            �����   +  >            �����   �   <   "         �����   �   =               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   ?            �����   +  B         	   ����      @      
      �����   �   A               ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   C            �����   +  D               ����                        ����                        ����                        ����                            +      #               �   E               �   +  J   !      	         �   F   #   
      �����   �   I   &         �����   �   K   0         �����   +  L   !         ����   �   G             �����   �   H               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   M            �����   +  N               ����                        ����                        ����                        ����                            +      +               �   O   *         �����   +  R         	   ����   �   P      
      �����   �   Q               ����                        ����                        ����                        ����                        ����                        ����                            +                     �   S   *         �����   +  X         	         �   T   #   
      �����   �   W               ����                        ����                     ����   �   U            �����   �   V               ����                        ����                        ����                        ����                        ����                        ����            "                +      +               �   Y            �����   +  ^         	         �   Z   +   
      �����   �   ]               ����                        ����                     ����   �   [            �����   �   \               ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   _   %         �����   +  `               ����                        ����                        ����                        ����                            +                     �   a            �����   +  f         	         W   b      
      ����X   �   e               ����                        ����                      ����      c            ����   W   d               ����                        ����                        ����                        ����                        ����                        ����                            +                     �   g            �����   +  j         	   ����   �   h      
      �����   �   i               ����                        ����                        ����                        ����                        ����                        ����                            +                     �   k               �   +  r         	         �   l      
      �����   �   q               �   '  s             ����(  +  z                  �   m            �����   �   p               ����                        ����                        �   �   t   *            �   '  w               ����                        ����                      �����   �   u   2         �����   �   v             �����   �   x            �����   '  y               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                   !   ����   �   n       "   #   �����   �   o               ����                        ����                        ����                        ����                        ����                        ����                            +      '         ����   �   {            �����   +  |               ����                        ����                        ����                        ����                            +                     �   }   *            �   +  �   $      	   ����      ~      
            �                �����   �   �            �����   +  �               ����                        ����                           �   �               �   �   �               ����                        ����                        ����                        ����            ,       !   ����   �   �       "   #   �����   �   �   '            �   �   �   %            �   �   �            �����   �   �   2         �����   �   �            �����   �   �            �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �               �   +  �               ����                        ����                  	      �   �   �   &   
         �   +  �            �����   �   �               �   �   �   *            �   �   �            �����   +  �            
   �   �   �   *         �����   �   �               ����                        ����                      �����   �   �             �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                     	   �   �   �            �����   �   �          !   �����   �   �   2   "   #   �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +      +               �   �            �����   +  �         	         �   �       
      �����   �   �               ����                        ����            $               �   �   1         �����   �   �               ����                        ����                     ����      �   $         ����   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �            �����   +  �         	   ����   �   �      
      �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �            �����   +  �         	         �   �      
         �   �   �               ����                        ����                     ����   �   �   1         �����   �   �   *         �����   �   �             �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �            �����   +  �         	         �   �   *   
         �   �   �               ����                        ����                      ����      �   !         ����   �   �   *         �����   �   �   *         �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �            �����   +  �         	         �   �      
      �����   �   �               ����                        ����                     ����   b   �            ����c   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �            �����   +  �   +      	   ����   ]   �      
      ����^   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �            �����   +  �   (      	   ����      �      
      ����   �   �               ����                        ����                        ����                        ����                        ����                        ����            #                +      "               �   �            �����   +  �   #      	   ����   �   �   	   
      �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +      +               �   �               �   +  �   '      	         �   �      
      �����   �   �            �����   �   �            �����   +  �                  �   �   '         �����   �   �               ����                        ����            !               �   �            �����   �   �               ����                        ����                           7   �               8   �   �               ����                        ����                        ����                        ����                        ����                        ����            '       !   ����      �      "   #         7   �             ����8   ;   �            ����<   �   �               ����                        ����                        ����                        ����                        ����                        ����            '   $   %   ����   $   �      &   '      %   7   �               ����                        ����            !   (   )   ����%   2   �       *   +   ����3   7   �               ����                        ����                        ����                        ����                            +                     �   �               �   +  �         	   ����   �   �   2   
      �����   �   �            �����   �   �            �����   +  �               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            "                +                     �   �            �����   +  �         	         �   �      
      �����   �   �               ����                        ����                     ����   W   �   $         ����X   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �            �����   +  �               ����                        ����                        ����                        ����                            +                     �   �               �   +  �         	         �   �      
      �����   �   �   2         �����   �   �            �����   +  �            ����   �   �   (         �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �   0            �   +  �               ����                        ����            !      	   �����   '  �       
      ����(  +  �               ����                        ����                        ����                        ����                            +                     �   �   0            �   +    )      	         �   �   2   
      �����   �                 �   &              ����'  +                   �   �            �����   �                  ����                        ����            "               �   �            �����   �   �               ����                        ����                     �����   �              �����   &                ����                        ����                        ����                        ����                        ����                        ����                     ����   �   �   )         �����   �   �               ����                        ����                        ����                        ����                        ����                        ����                            +      '         ����   �              �����   +                ����                        ����                        ����                        ����                            +                     �   	           �����   +    *      	         }   
     
         ~   �                 ����                        ����            '                             ����   }              ����~   �              �����   �     1         ����        *         ����                    ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      +         ����   �              �����   +                ����                        ����                        ����                        ����            #                +                     �              �����   +          	   ����   �     #   
      �����   �                 ����                        ����                        ����                        ����                        ����                        ����                            +                     �              �����   +  "  '      	         �     2   
      �����   �   !              ����                        ����                     ����   �                 �   �                 ����                        ����                        ����                        ����                      �����   �              	   �   �                 ����                        ����            2         �����   �              �����   �                  ����                        ����                        ����                        ����                            +               ����   V   #              W   +  $              ����                        ����                  	   ����W   �   %  *   
      �����   +  &              ����                        ����                        ����                        ����            #                +                     �   '  !            �   +  *  *      	   ����   �   (     
      �����   �   )           �����   $  +  (         ����%  +  ,              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      )         ����   �   -  *         �����   +  .              ����                        ����                        ����                        ����                            +      +         ����   �   /           �����   +  0              ����                        ����                        ����                        ����            /                +               ����   �   1  /         �����   +  2              ����                        ����                        ����                        ����                            +                     �   3  ,         �����   +  8  '      	   ����      4  !   
            �   5              ����                        ����                        ����                        ����                     ����   �   6            �����   �   7              ����                        ����                        ����                        ����                            +      '               �   9  0         �����   +  <        	   ����   �   :  '   
      �����   �   ;              ����                        ����                        ����                        ����                        ����                        ����            #                +      #         ����   �   =  %            �   +  >              ����                        ����                   	   �����   �   ?  0   
         �   +  @              ����                        ����            +            �   '  A            ����(  +  D  0         �����   �   B  *         �����   '  C              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   E           �����   +  F              ����                        ����                        ����                        ����                            +               ����   �   G           �����   +  H              ����                        ����                        ����                        ����                            +               ����   �   I           �����   +  J              ����                        ����                        ����                        ����                            +      '         ����   �   K  *         �����   +  L              ����                        ����                        ����                        ����                            +                     �   M           �����   +  P        	   ����   �   N     
      �����   �   O              ����                        ����                        ����                        ����                        ����                        ����            #                +      #         ����   �   Q  !            �   +  R              ����                        ����                  	      �   !  S  #   
      ����"  +  V            �����   �   T  )         �����   !  U              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   W           �����   +  Z        	   ����   �   X  2   
      �����   �   Y              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   [  *         �����   +  b  ,      	         �   \     
      �����   �   a              ����                        ����            ,               �   ]            �����   �   `              ����                        ����                     ����   �   ^           �����   �   _              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   c           �����   +  f        	   ����      d     
      ����	   �   e              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   g              �   +  h              ����                        ����                  	   �����   �   i  *   
         �   +  j              ����                        ����                     �����   &  k            ����'  +  l              ����                        ����                        ����                        ����                            +                     �   m           �����   +  |        	            n     
            �   q              ����                        ����                     ����      o            ����      p           ����   \   r              ]   �   s              ����                        ����                        ����                        ����                        ����                        ����                        ]   �   t           �����   �   {              ]   f   u  0            g   �   x              ����                        ����                    !   ����]   `   v  2   "   #   ����a   f   w           ����g   �   y  0         �����   �   z              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      $               �   }  #         �����   +  �        	   ����   �   ~     
      �����   �                 ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	         �   �      
      �����   �   �              ����                        ����                           �   �           �����   �   �              ����                        ����            %         ����   �   �           �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �  0   
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �              �   +  �        	         �   �     
      �����   �   �           �����     �           ����  +  �           ����   �   �           �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      '               �   �           �����   +  �  0      	         �   �     
      �����   �   �              ����                        ����            /               �   �  1         �����   �   �              ����                        ����            '         ����   �   �  1         �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����      �     
      ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �  *         �����   +  �              ����                        ����                        ����                        ����                            +                     �   �  !            �   +  �        	   ����   j   �     
      ����k   �   �           �����   '  �            ����(  +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            #                +      #         ����   �   �           �����   +  �              ����                        ����                        ����                        ����                            +                     �   �  *            �   +  �        	         ^   �     
         _   �   �              �   �   �  *         �����   +  �                 
   �                 ^   �         !      _   �   �      "   #   �����   �   �           �����   �   �  2         �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                      ����      �            ����   
   �           	      X   �  2         ����Y   ^   �     D   E         -   �     F   G   ����.   X   �              ����                        ����                        ����                        ����                        ����                        ����               $   %   
   _   �   �  '   &   '   
   �   �   �              ����                        ����               ,   -   ����_   t   �  	   .   /       u   �   �     (   )   �����   �   �  %   *   +   !   �   �   �              ����                        ����                0   1   �����   �   �     2   3   �����   �   �              ����                        ����            	   4   5   %   u   �   �     6   7   �����   �   �              ����                        ����                        ����                        ����               8   9   .   u   �   �      :   ;   �����   �   �              ����                        ����            	   <   =   ����u   {   �  *   >   ?   4   |   �   �              ����                        ����                        ����                        ����                @   A   ����|   �   �  	   B   C   �����   �   �              ����                        ����                        ����                        ����            %   H   I   ����      �     J   K         -   �              ����                        ����                        ����                        ����            *   L   M   ����   %   �     N   O   ����&   -   �              ����                        ����                        ����                        ����                            +                     �   �  *         �����   +  �        	   ����   �   �     
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �           �����   +  �              ����                        ����                        ����                        ����                            +                     �   �  ,         �����   +  �        	         �   �     
      �����   �   �              ����                        ����                      ����      �           ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �  !   
         �   �   �              ����                        ����                        ����                        ����            %         �����   �   �  !         �����   �   �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �     
         �   �   �              ����                        ����                        ����                        ����                        �   �   �              �   �   �            �����   �   �           �����   �   �           �����   �   �            �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            #                +      /               �   �  !         �����   +  �  #      	   ����   �   �      
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �  *         �����   +  �        	         �   �  1   
         �   �   �              ����                        ����                     ����   �   �           �����   �   �           �����   �   �              �   �   �              ����                        ����            1         �����   �   �            �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +           	         �   �     
      �����   �   �              ����                        ����                     ����   �   �           �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �     +            �   +                ����                        ����                  	   �����   '        
      ����(  +                ����                        ����                        ����                        ����                            +      '               �              �����   +          	   ����   �        
      �����   �                 ����                        ����                        ����                        ����                        ����                        ����                            +      $               �   	  !            �   +    $         ����   �   
           �����   �           	   �����   '        
      ����(  +                ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �     (         �����   +          	         �        
      �����   �                 ����                        ����                     ����   l              ����m   �                 ����                        ����                        ����                        ����                        ����                        ����            )                +      ,               �     )         �����   +    +      	         �        
      �����   �                 ����                        ����                     ����   �     2         �����   �                 ����                        ����                        ����                        ����                        ����                        ����                            +      	         ����   �     )         �����   +                ����                        ����                        ����                        ����                            +                     �                 �   +  6        	         {        
         |   �   #      0   1   �����   �   7  %   2   3   �����   +  8     4   5         r        6   7   ����s   {   "              |   �   $  1            �   �   +  '   $   %   
   |   �   %     &   '   �����   �   *  1         �����   �   ,              �   �   -              ����                        ����                        �   �   .              �   �   3              �   �   /           �����   �   2            �����   �   4  #         �����   �   5              ����                        ����                        ����                        ����            1       !   �����   �   0      "   #   �����   �   1              ����                        ����                        ����                        ����                        ����                        ����               (   )      |   �   &  2   *   +   �����   �   )              ����                        ����               ,   -   ����|   �   '     .   /   �����   �   (              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            +   8   9   ����   c         :   ;   ����d   r   !              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   9           �����   +  <        	   ����   �   :     
      �����   �   ;              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   =           �����   +  @        	   ����   y   >     
      ����z   �   ?              ����                        ����                        ����                        ����                        ����                        ����                            +      $               [   A              \   +  D  $         ����   W   B            ����X   [   C  '      	      \   �   E  *   
         �   +  H  '         ����\   �   F           �����   �   G           �����   �   I           �����   +  J              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   K              �   +  L              ����                        ����                  	   �����   %  M  2   
      ����&  +  N              ����                        ����                        ����                        ����                            +      0               �   O  *         �����   +  T  .      	         �   P  (   
      �����   �   S              ����                        ����            '         ����   �   Q            �����   �   R              ����                        ����                        ����                        ����                        ����                        ����            #                +      #               �   U  #         �����   +  X  *      	   ����   j   V     
      ����k   �   W              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   Y           �����   +  \        	   ����   w   Z     
      ����x   �   [              ����                        ����                        ����                        ����                        ����                        ����                            +      $               �   ]  #         �����   +  b        	   ����   =   ^     
         >   �   _              ����                        ����                        ����                        ����            1         ����>   �   `           �����   �   a              ����                        ����                        ����                        ����                            +                     �   c           �����   +  f        	   ����   n   d     
      ����o   �   e              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   g           �����   +  h              ����                        ����                        ����                        ����                            +                     �   i           �����   +  t  $      	            j  +   
            �   o              ����                        ����                              k  1         ����      n                 �   p            �����   �   s  1         ����   }   q  2         ����~   �   r              ����                        ����                        ����                        ����                        ����                        ����                      ����      l           ����      m              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   u              �   +  x        	   ����   �   v     
      �����   �   w           �����   �   y  )         �����   +  z              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            #                +                     �   {  #         �����   +  �        	         �   |  1   
      �����   �   �              ����                        ����                     ����   +   }  *            ,   �   ~              ����                        ����                        ����                        ����            $         ����,   ]     *         	   ^   �   �              ����                        ����                     ����^   x   �              y   �   �              ����                        ����            #         ����y   �   �  *         �����   �   �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	         �   �      
      �����   �   �              ����                        ����            2         ����   e   �           ����f   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �  0            �   +  �        	   ����   `   �     
         a   �   �              �   &  �            ����'  +  �              ����                        ����                     ����a   �   �              �   �   �              ����                        ����                     �����   �   �            �����   �   �           �����   !  �            ����"  &  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �  !         �����   +  �  1      	   ����      �  '   
      ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +      !               �   �  *         �����   +  �        	   ����      �     
             �   �              ����                        ����                        ����                        ����            2         ����    �   �  2         �����   �   �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	         �   �      
      �����   �   �              ����                        ����                     ����   �   �           �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �  0         �����   +  �        	   ����   �   �      
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            )                +      +               �   �  )         �����   +  �  +      	   ����   �   �  2   
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            #                +      #         ����   �   �              �   +  �              ����                        ����                  	   �����   �   �  #   
      �����   +  �              ����                        ����                        ����                        ����                            +                     �   �  ,         �����   +  �  '      	   ����   �   �     
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            )                +      )         ����   �   �           �����   +  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����      �     
            �   �              ����                        ����                        ����                        ����                     ����   �   �              �   �   �              ����                        ����                     �����   �   �           �����   �   �              ����                        ����                        ����                        ����                            +               ����   �   �  *         �����   +  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �      
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �  1   
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +      *               �   �              �   +  �         	   ����      �  *   
      ����   �   �           �����   �   �           �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �  *         �����   +  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	         �   �     
      �����   �   �              ����                        ����            $               �   �           �����   �   �              ����                        ����            $         ����   �   �  $            �   �   �              ����                        ����                        ����                        ����            1         �����   �   �  $            �   �   �              ����                        ����                      �����   �   �  $         �����   �   �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �         	   ����      �  $   
      ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +      ,               �   �           �����   +  �        	         (   �     
      ����)   �   �              ����                        ����            ,         ����      �  ,         ����   (   �              ����                        ����                        ����                        ����                        ����                        ����            #                +      *               �   �  #         �����   +  �  #      	   ����   �   �      
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            *                +      *         ����   K   �           ����L   +  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	         j   �      
         k   �   �              ����                        ����            *         ����   	   �           ����
   j   �           ����k   �   �  -         �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            *                +      *         ����   g   �              h   +  �              ����                        ����                  	      h   �   �     
      �����   +  �  (         ����h   �   �           �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +      	               �   �           �����   +    '      	   ����   �         
      �����   �                 ����                        ����                        ����                        ����                        ����                        ����            *                +                     �     *         �����   +    +      	         w        
      ����x   �                 ����                        ����            +               p     *         ����q   w                 ����                        ����            $               h     *         ����i   p                 ����                        ����                           a                 b   h   
              ����                        ����            $         ����   ]               ����^   a   	            ����b   d               ����e   h                 ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �                 �   +  ,        	         9        
         :   �              �����     -                +  .      $   %   ����           &   '   ����   9     ,            :   �              �����   �   +              ����                        ����                      ����     /           ����!  +  0              ����                        ����                        ����                        ����            ,         
   :   l     ,         
   m   �                 ����                        ����                     ����:   @     $            A   l        ,   -      m   �        .   /      �   �   &              ����                        ����                   !      A   R     ,   "   #   ����S   l     1   (   )   ����A   F     $   *   +   ����G   R                 ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����               0   1      m   �          2   3   �����   �   %  1   4   5   �����   �   '  *   6   7      �   �   (  "   8   9   ,   m   �   !      :   ;   �����   �   $              ����                        ����                        ����                        ����                @   A   �����   �   )      B   C   �����   �   *     <   =   ����m   �   "      >   ?   �����   �   #              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      '               �   1           �����   +  4  *      	   ����   �   2  2   
      �����   �   3              ����                        ����                        ����                        ����                        ����                        ����                            +      '               �   5  *         �����   +  :        	         �   6     
      �����   �   9              ����                        ����                      ����      7           ����   �   8              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   ;  #         �����   +  <              ����                        ����                        ����                        ����                            +               ����   �   =  !         �����   +  >              ����                        ����                        ����                        ����                            +                     `   ?           ����a   +  B        	   ����   0   @  %   
      ����1   `   A              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   C           �����   +  F        	   ����   �   D     
      �����   �   E              ����                        ����                        ����                        ����                        ����                        ����                            +      +               �   G           �����   +  J  '      	   ����   �   H  2   
      �����   �   I              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   K  0         �����   +  L              ����                        ����                        ����                        ����                            +      ,               |   M           ����}   +  P  ,      	   ����   Y   N  +   
      ����Z   |   O              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   Q           �����   +  T        	   ����   	   R  '   
      ����
   �   S              ����                        ����                        ����                        ����                        ����                        ����                            +      "         ����   �   U           �����   +  V              ����                        ����                        ����                        ����            *                +                     p   W           ����q   +  Z        	   ����   `   X     
      ����a   p   Y              ����                        ����                        ����                        ����                        ����                        ����                            +      '               |   [  #         ����}   +  ^  '      	   ����   t   \  1   
      ����u   |   ]              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   _           �����   +  `              ����                        ����                        ����                        ����                            +                     �   a  (            �   +  f                 �   b           �����   �   e         	   �����   �   g  (   
      �����   +  h              ����                        ����                        ����                        ����            -         ����   �   c            �����   �   d              ����                        ����                        ����                        ����                        ����                        ����            "                +      "               �   i  "         �����   +  l  2      	   ����   �   j     
      �����   �   k              ����                        ����                        ����                        ����                        ����                        ����            "                +                     �   m           �����   +  r        	   ����   	   n     
         
   �   o              ����                        ����                        ����                        ����                     ����
   E   p           ����F   �   q              ����                        ����                        ����                        ����                            +      *         ����   �   s           �����   +  t              ����                        ����                        ����                        ����                            +      !         ����   �   u           �����   +  v              ����                        ����                        ����                        ����                            +               ����   
   w                 +  x              ����                        ����                  	         �   y     
         �   +  |  0         ����   �   z           �����   �   {  #         �����     }  )         ����  +  ~              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �     0         �����   +  �              ����                        ����                        ����                        ����            *                +      '         ����   m   �              n   +  �              ����                        ����                  	   ����n   �   �  *   
      �����   +  �              ����                        ����                        ����                        ����                            +               ����   �   �           �����   +  �              ����                        ����                        ����                        ����                            +                     �   �  *            �   +  �  %      	   ����      �     
      ����   �   �           �����   �   �           �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �  ,   
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            )                +      )         ����   �   �  )            �   +  �              ����                        ����                   	   �����   �   �  )   
         �   +  �              ����                        ����            )            �   �   �  )         �����   +  �           �����   �   �            �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   P   �     
         Q   �   �              ����                        ����                        ����                        ����                     ����Q   n   �              o   �   �              ����                        ����            1         ����o   x   �  #         ����y   �   �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �         	   ����      �     
            �   �              ����                        ����                        ����                        ����                     ����   t   �           ����u   �   �              ����                        ����                        ����                        ����                            +      1               �   �              �   +  �  1      	   ����   l   �  1   
      ����m   �   �  1         �����   �   �           �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            *                +      '               �   �  *         �����   +  �  *      	         �   �  *   
         �   �   �              ����                        ����            *         ����   d   �  '            e   �   �  1         �����   �   �              �   �   �              ����                        ����            *         ����e   �   �  *         �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            '         �����   �   �           �����   �   �              ����                        ����                        ����                        ����                            +      ,               �   �  0            �   +  �  ,      	   ����   Q   �  ,   
      ����R   �   �  *         �����   $  �  .            %  +  �              ����                        ����                        ����                        ����                        ����                        ����                      ����%  '  �            ����(  +  �              ����                        ����                        ����                        ����            *                +      *         ����   �   �           �����   +  �              ����                        ����                        ����                        ����            #                +      #               �   �  #         �����   +  �  ,      	   ����   d   �  /   
      ����e   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �              �   +  �  #               �   �  -         �����   �   �        	   �����   �   �     
         �   +  �              ����                        ����                        �   �   �  $         �����   +  �           
   �   �   �  #         �����   �   �              ����                        ����                      �����   �   �            �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            #         ����   t   �  #         ����u   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +      $               �   �           �����   +  �        	         d   �  $   
      ����e   �   �              ����                        ����                     ����   ^   �  2         ����_   d   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �              �   +  �              ����                        ����                  	   �����   &  �      
      ����'  +  �              ����                        ����                        ����                        ����                             +                ����      �                 +  �              ����                        ����                  	         �   �     
         �   +  �           ����   "   �            ����#   �   �           �����   $  �              %  +  �              ����                        ����                        ����                        ����                        ����                        ����                      ����%  '  �            ����(  +  �              ����                        ����                        ����                        ����            '                +                       �                +  �        	         �   �  *   
      �����     �            ����    �                +  �                 �   �            �����   �   �              ����                        ����                        ����                        ����            '   $   %   ����     �     &   '   ����!  +  �                 �   �  '            �   �   �              ����                        ����                           
   �           ����   �   �          !   �����   �   �     "   #   �����   �   �            ����      �  2         ����   
   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �     
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �  $            �   +           	   ����            
      ����   �     *         �����   �     $         �����   +                ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            *                +                ����   �              �����   +                ����                        ����                        ����                        ����                            +                     �              �����   +          	         a        
      ����b   �                 ����                        ����                     ����   X   	  $         ����Y   a   
              ����                        ����                        ����                        ����                        ����                        ����                            +      $         ����   �              �����   +                ����                        ����                        ����                        ����                            +               ����   �              �����   +                ����                        ����                        ����                        ����                            +      $               �              �����   +    #      	   ����   �     $   
      �����   �                 ����                        ����                        ����                        ����                        ����                        ����            )                +      )               �     !            �   +    )               �               �����   �     )      	   �����   &        
      ����'  +                 ����                        ����                        ����                        ����                            �     )            �   �                 ����                        ����                      ����        )         ����   �     )         �����   �               �����   �                 ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   !           �����   +  $        	   ����   �   "      
      �����   �   #              ����                        ����                        ����                        ����                        ����                        ����            *                +                     i   %  *         ����j   +  *  *      	         b   &  *   
      ����c   i   )              ����                        ����                     ����      '  *         ����   b   (              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   +           �����   +  .        	   ����   �   ,  +   
      �����   �   -              ����                        ����                        ����                        ����                        ����                        ����            )                +      )         ����   �   /  )         �����   +  0              ����                        ����                        ����                        ����            #                +      #               �   1  #         �����   +  8        	         �   2  2   
      �����   �   7              ����                        ����                           �   3            �����   �   6              ����                        ����                     ����   i   4           ����j   �   5              ����                        ����                        ����                        ����                        ����                        ����            +                +                     �   9              �   +  F  +      	         �   :  +   
      �����   �   E           �����   �   G           �����   +  H                 �   ;           �����   �   D              ����                        ����                        ����                        ����                        ����                        ����                     ����   i   <               j   �   =              ����                        ����                        ����                        ����            ,            j   �   >              �   �   A            ����j   l   ?           ����m   �   @         !   �����   �   B  '   "   #   �����   �   C              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +                     �   I  ,         �����   +  P        	         �   J     
      �����   �   O              ����                        ����            $               �   K            �����   �   N              ����                        ����                     ����      L  $         ����    �   M              ����                        ����                        ����                        ����                        ����                        ����                            +                        Q           ����  +  T  '      	   ����   �   R      
      �����      S              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   U              �   +  ^        	         �   V     
         �   �   [           �����   �   _           �����   +  `           ����   �   W  *            �   �   X           �����   �   \           �����   �   ]              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                      �����   �   Y  )         �����   �   Z              ����                        ����                        ����                        ����                            +      ,         ����   �   a           �����   +  b              ����                        ����                        ����                        ����            $                +                ����      c  $               +  d              ����                        ����                  	   ����      e  $   
            +  f              ����                        ����            $         ����   (   g  %            )   +  h              ����                        ����            %         ����)   �   i  '            �   +  j              ����                        ����                        �   #  k  '         ����$  +  n  '         �����   �   l  %         �����   #  m              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   o  #         �����   +  t  !      	         �   p  $   
      �����   �   s              ����                        ����            !         ����   -   q           ����.   �   r              ����                        ����                        ����                        ����                        ����                        ����            *                +      %         ����   d   u           ����e   +  v              ����                        ����                        ����                        ����                            +      '               �   w  #         �����   +  z        	   ����   �   x  '   
      �����   �   y              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   {           �����   +  ~        	   ����   �   |     
      �����   �   }              ����                        ����                        ����                        ����                        ����                        ����            "                +               ����   �     "         �����   +  �              ����                        ����                        ����                        ����            1                +               ����   +   �              ,   +  �              ����                        ����                  	   ����,   �   �  2   
      �����   +  �              ����                        ����                        ����                        ����                            +               ����   a   �  %         ����b   +  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   �   �      
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����      �     
      ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	         �   �     
      �����   �   �              ����                        ����            (         ����   �   �  ,         �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �  )            �   +  �        	         �   �     
      �����   �   �            �����   �   �  )         �����   +  �            ����      �           ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            '                +      %         ����     �  '         ����  +  �              ����                        ����                        ����                        ����            '                +                       �  '         ����  +  �  )      	   ����   
   �  !   
      ����     �              ����                        ����                        ����                        ����                        ����                        ����                            +      .               �   �              �   +  �  .      	   ����   �   �      
      �����   �   �           �����   �   �           �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            .                +      -               �   �           �����   +  �        	         �   �  $   
      �����   �   �              ����                        ����            *               -   �           ����.   �   �              ����                        ����                     ����   '   �  2         ����(   -   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �              �   +  �              ����                        ����                   	   �����   �   �     
      �����   +  �              ����                        ����                        ����                        ����            *                +                      "   �              #   +  �  1         ����      �  *         ����   "   �        	   ����#   �   �     
      �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            +                +      0         ����   �   �           �����   +  �              ����                        ����                        ����                        ����            *                +                        �  *         ����   +  �         	   ����      �  *   
      ����      �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �              �   +  �           ����      �                 �   �        	   �����     �  '   
           +  �              ����                        ����                     ����    �  '         ����  +  �              ����                        ����                        ����                        ����                        ����                        ����            ,               �   �            �����   �   �  ,         ����   !   �              "   �   �              ����                        ����                        ����                        ����            ,         ����"   �   �           �����   �   �              ����                        ����                        ����                        ����                            +               ����   �   �  *         �����   +  �              ����                        ����                        ����                        ����            "                +      -               �   �  "         �����   +  �         	         �   �  -   
      �����   �   �              ����                        ����                      ����      �            ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     u   �              v   +  �         	   ����      �     
      ����   u   �            ����v   z   �              {   +  �              ����                        ����                        ����                        ����                        ����                        ����                        {   �   �              �   +  �           ����{   �   �           �����   �   �  *         �����   �   �  *         �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �  #            �   +  �              ����                        ����                   	   �����   �   �     
      �����   +  �              ����                        ����                        ����                        ����            *                +      *         ����   q   �  *            r   +  �              ����                        ����            2      	   ����r   w   �  *   
      ����x   +  �              ����                        ����                        ����                        ����                            +                     �   �  ,            �   +  �           ����      �  *         ����   �   �  /      	   �����   �   �  ,   
      �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      "               �   �           �����   +  �        	   ����   �   �     
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �              �   +  �        	   ����      �     
      ����	   �   �              �   �   �              �   +  �              ����                        ����                        ����                        ����                     �����   �   �            �����   �   �           �����   �   �  )         �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +               ����     �  *              +                 ����                        ����            #      	   ����      *   
      ����  +                ����                        ����                        ����                        ����            '                +                         '         ����  +    '      	         �     $   
         �                   ����                        ����            ,         ����   p     '         ����q   �               �����   �                 �     	              ����                        ����                     �����     
            ����	                  ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            (                +               ����   M                 N   +                ����                        ����                  	   ����N           
      ����  +                ����                        ����                        ����                        ����                            +                     �                 �   +           	   ����           
      ����   �     /         �����   �              �����   +                ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      *               �     !         �����   +          	   ����   [     *   
      ����\   �                 ����                        ����                        ����                        ����                        ����                        ����            *                +      $               c     ,            d   +           	   ����        *   
      ����   c     '         ����d   o              ����p   +                 ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            +                +      +               �   !  *         �����   +  &        	         �   "  +   
      �����   �   %              ����                        ����                     ����   �   #            �����   �   $              ����                        ����                        ����                        ����                        ����                        ����            '                +      )         ����   �   '  ,            �   +  (              ����                        ����            '      	   �����     )  ,   
      ����  +  *              ����                        ����                        ����                        ����                            +               ����     +           ����  +  ,              ����                        ����                        ����                        ����                            +               ����   �   -           �����   +  .              ����                        ����                        ����                        ����            '                +      '         ����     /  '              +  0              ����                        ����            #      	   ����    1  '   
      ����  +  2              ����                        ����                        ����                        ����                            +      !         ����   �   3  $         �����   +  4              ����                        ����                        ����                        ����                             +                ����     5                 +  6              ����                        ����            #      	   ����    7  1   
      ����  +  8              ����                        ����                        ����                        ����                            +      )         ����      9                 +  :              ����                        ����                  	         �   ;     
      �����   +  F                 z   <           ����{   �   E              ����                        ����            !               @   =           ����A   z   D              ����                        ����            !               :   >  2         ����;   @   C              ����                        ����            +               6   ?            ����7   :   B              ����                        ����                     ����   *   @  )         ����+   6   A              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   G  !         �����   +  H              ����                        ����                        ����                        ����                            +      '         ����   �   I  *            �   +  J              ����                        ����            2      	   �����   �   K  *   
      �����   +  L              ����                        ����                        ����                        ����                            +                     �   M              �   +  X  ,               �   N           �����   �   W        	   �����   �   Y     
      �����   +  Z              ����                        ����                        ����                        ����            ,               e   O              f   �   T              ����                        ����                     ����      P                 e   Q           ����f   �   U  1         �����   �   V              ����                        ����                        ����                        ����                        ����                        ����                     ����   ^   R  ,         ����_   e   S              ����                        ����                        ����                        ����                            +                     �   [           �����   +  ^        	   ����   �   \      
      �����   �   ]              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   _           �����   +  `              ����                        ����                        ����                        ����            0                +      0               $  a  '         ����%  +  d        	   ����   �   b  0   
      �����   $  c              ����                        ����                        ����                        ����                        ����                        ����                            +      *         ����      e  0               +  f              ����                        ����            0      	         $  g      
         %  +  t  0               �   h  0         �����   $  s            ����%  '  u            ����(  +  v  0               �   i              �   �   p              ����                        ����                        ����                        ����                        ����                        ����                           �   j            �����   �   o  0         �����   �   q           �����   �   r              ����                        ����                        ����                        ����                   !   ����   a   k     "   #      b   �   l              ����                        ����                        ����                        ����                $   %   ����b   e   m     &   '   ����f   �   n              ����                        ����                        ����                        ����                            +      0               y   w           ����z   +  z  +      	   ����   s   x  2   
      ����t   y   y              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   t   {              u   +  |              ����                        ����            ,      	   ����u   �   }     
      �����   +  ~              ����                        ����                        ����                        ����                            +      *         ����   �              �����   +  �              ����                        ����                        ����                        ����                            +                     	  �           ����
  +  �        	   ����   (   �  .   
         )   	  �              ����                        ����                        ����                        ����            '         ����)   �   �           �����   	  �              ����                        ����                        ����                        ����            +                +      +               �   �              �   +  �  +         ����   �   �              �   �   �  2      	   �����   �   �  +   
      �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                     �����   �   �  +         �����   �   �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����      �  '   
      ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �              �   +  �              ����                        ����                  	   �����     �     
      ����  +  �              ����                        ����                        ����                        ����                            +                     -   �              .   +  �        	   ����      �  &   
            -   �  1            .   '  �            ����(  +  �              ����                        ����            #               &   �  &         ����'   -   �           ����       �  2         ����!   &   �              ����                        ����                        ����                        ����                        ����                        ����                     ����.   �   �              �   '  �              ����                        ����                        ����                        ����            ,            �   �   �           ����   '  �         !   �����   �   �     "   #      �   �   �              ����                        ����                        ����                        ����               $   %   �����   �   �     &   '   �����   �   �              ����                        ����                        ����                        ����                            +      +         ����   d   �  '            e   +  �              ����                        ����                  	      e   	  �     
      ����
  +  �           ����e   �   �           �����   	  �              ����                        ����                        ����                        ����                        ����                        ����                            +      )               l   �           ����m   +  �        	   ����   S   �  )   
      ����T   l   �              ����                        ����                        ����                        ����                        ����                        ����                            +                     $  �  1         ����%  +  �        	   ����   a   �  #   
         b   $  �              ����                        ����                        ����                        ����                     ����b   �   �  #         �����   $  �              ����                        ����                        ����                        ����                            +                     '  �            ����(  +  �        	           �     
      ����  '  �              ����                        ����            )         ����   �   �  $            �     �              ����                        ����                        ����                        ����            #         �����   �   �  $         �����     �              ����                        ����                        ����                        ����            )                +               ����   �   �  )         �����   +  �              ����                        ����                        ����                        ����            '                +      '         ����   �   �  ,            �   +  �              ����                        ����            1      	   �����   �   �     
      �����   +  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �  ,      	         n   �     
      ����o   �   �              ����                        ����            ,         ����   8   �           ����9   n   �              ����                        ����                        ����                        ����                        ����                        ����            '                +      &               �   �  ,            �   +  �  '      	   ����   j   �  $   
      ����k   �   �  '         �����   �   �           �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            +      '               �   �  0            �   +  �           ����   �   �           �����   �   �        	   �����   '  �      
      ����(  +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            1                +               ����      �  *            	   +  �              ����                        ����            )      	      	   `   �  1   
         a   +  �              	   W   �  1         ����X   `   �              a   �   �  *         �����   +  �  *         ����	   S   �            ����T   W   �              ����                        ����                        ����                        ����                        ����                        ����            *         ����a   �   �  )         
   �   �   �              ����                        ����                        ����                        ����            *         �����   �   �  )         �����   �   �              ����                        ����                        ����                        ����                             +      ,               �   �            �����   +  �        	   ����   X   �     
         Y   �   �              ����                        ����                        ����                        ����                     ����Y   �   �           �����   �   �              ����                        ����                        ����                        ����            +                +      +               �   �           �����   +  �        	         �   �     
      �����   �   �              ����                        ����            *         ����   �   �  *            �   �   �              ����                        ����                        ����                        ����            '         	   �   �   �  *         �����   �   �           �����   �   �  ,         �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            	                +      $                 �                +  �  $      	   ����      �     
              �           ����  &  �            ����'  +                 ����                        ����            $         ����   j   �  	            k     �              ����                        ����            2         ����k   p   �           ����q     �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            #                +      #         ����   �     #         �����   +                ����                        ����                        ����                        ����                            +               ����   �                 �   +                ����                        ����            !      	   �����   �        
      �����   +                ����                        ����                        ����                        ����                            +                     �              �����   +          	         �     #   
         �   �                 ����                        ����                     ����   �   	            �����   �   
            �����   �              �����   �                 ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            %                +      	         ����   �     %         �����   +                ����                        ����                        ����                        ����                            +                     �     .            �   +                   r                 s   �           	      �       .   
      ����  +    2         �����                ����                  ����                        ����                        ����                        ����                        ����                        ����                     ����   S              ����T   r     0         ����s   �              �����   �                 ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            *                +                      m     *         ����n   +  $  (      	         b         
      ����c   m   #              ����                        ����            2               ]               ����^   b   "              ����                        ����            '         ����   X                ����Y   ]   !              ����                        ����                        ����                        ����                        ����                        ����            '                +      !                 %  '         ����  +  ,        	           &  2   
      ����    +              ����                        ����            '         ����      '                   (              ����                        ����                        ����                        ����                     ����   �   )           �����     *              ����                        ����                        ����                        ����                            +      ,         ����      -           ����   +  .              ����                        ����                        ����                        ����            /                +      1         ����   �   /  /         �����   +  0              ����                        ����                        ����                        ����            &                +      &               �   1  &         �����   +  8  &      	         �   2     
         �   �   5              ����                        ����            &         ����   �   3  &         �����   �   4            �����   �   6            �����   �   7              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                             +               ����      9           ����   +  :              ����                        ����                        ����                        ����                            +               ����   i   ;  '            j   +  <              ����                        ����                  	   ����j     =     
      ����  +  >              ����                        ����                        ����                        ����                            +      (         ����      ?                 +  @              ����                        ����                  	   ����   Y   A  *   
      ����Z   +  B              ����                        ����                        ����                        ����            *                +                     l   C  *         ����m   +  F        	   ����   Z   D     
      ����[   l   E              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   G           �����   +  H              ����                        ����                        ����                        ����                            +               ����   G   I              H   +  J              ����                        ����            $      	   ����H   P   K     
      ����Q   +  L              ����                        ����                        ����                        ����            '                +      '         ����     M  (         ����  +  N              ����                        ����                        ����                        ����            #                +                     �   O  #         �����   +  R  #      	   ����   �   P      
      �����   �   Q              ����                        ����                        ����                        ����                        ����                        ����            0                +      0               �   S  0            �   +  X  +               �   T           �����   �   W        	   �����   	  Y  0   
      ����
  +  Z              ����                        ����                        ����                        ����            1         ����   �   U  +         �����   �   V              ����                        ����                        ����                        ����                        ����                        ����            !                +      !         ����   '  [            ����(  +  \              ����                        ����                        ����                        ����            '                +      !         ����     ]  '         ����  +  ^              ����                        ����                        ����                        ����                            +                     \   _           ����]   +  b         	   ����      `     
      ����   \   a              ����                        ����                        ����                        ����                        ����                        ����            '                +      '               $  c           ����%  +  f  0      	   ����   �   d  ,   
      �����   $  e              ����                        ����                        ����                        ����                        ����                        ����            	                +      	         ����   �   g           �����   +  h              ����                        ����                        ����                        ����            %                +      %               �   i  %         �����   +  n         	   ����      j  1   
            �   k              ����                        ����                        ����                        ����            1         ����   u   l  %         ����v   �   m              ����                        ����                        ����                        ����            +                +      '               �   o           �����   +  t        	         �   p     
      �����   �   s              ����                        ����            +         ����   �   q  '         �����   �   r              ����                        ����                        ����                        ����                        ����                        ����            *                +      *               y   u  *         ����z   +  z  '      	         d   v  )   
      ����e   y   y              ����                        ����            '         ����   `   w            ����a   d   x              ����                        ����                        ����                        ����                        ����                        ����                            +                        {           ����   +  ~        	   ����      |     
      ����      }              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �     *            �   +  �              ����                        ����            *      	   �����   �   �     
      �����   +  �              ����                        ����                        ����                        ����            *                +      !               j   �  *            k   +  �  !      	   ����   d   �  2   
      ����e   j   �            ����k   m   �              n   +  �              ����                        ����                        ����                        ����                        ����                        ����            *         ����n   {   �  )            |   +  �              ����                        ����            )         ����|   �   �  *         �����   +  �              ����                        ����                        ����                        ����            !                +      !               '  �            ����(  +  �        	   ����   #  �      
      ����$  '  �              ����                        ����                        ����                        ����                        ����                        ����                             +                      �   �              �   +  �  *         ����   X   �           ����Y   �   �  )      	   �����   �   �      
      �����   +  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            !                +                     "  �  2         ����#  +  �        	         �   �     
      �����   "  �              ����                        ����            !                  �                 �   �              ����                        ����            '       !   ����      �      "   #   ����	      �  !         	      z   �           	   {   �   �                 j   �              k   z   �  !   $   %   ����{   �   �  !   &   '   �����   �   �           ����   R   �           ����S   j   �           ����k   s   �  !         ����t   z   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                             +                ����      �                 +  �              ����                        ����            +      	   ����   u   �     
      ����v   +  �              ����                        ����                        ����                        ����            (                +               ����      �                 +  �              ����                        ����                  	            �     
      ����   +  �            ����      �  (         ����      �              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����   q   �     
      ����r   �   �              ����                        ����                        ����                        ����                        ����                        ����            '                +      '                 �  '         ����  +  �        	   ����   C   �     
      ����D     �              ����                        ����                        ����                        ����                        ����                        ����            !                +      !         ����   9   �              :   +  �              ����                        ����                  	      :   �   �     
      �����   +  �           ����:   �   �           �����   �   �              ����                        ����                        ����                        ����                        ����                        ����            !                +      *         ����   �   �           �����   +  �              ����                        ����                        ����                        ����                            +               ����     �                +  �              ����                        ����                   	   ����    �     
           +  �              ����                        ����                     ����  "  �           ����#  +  �              ����                        ����                        ����                        ����                            +                        �           ����   +  �         	   ����      �  #   
      ����      �              ����                        ����                        ����                        ����                        ����                        ����            *                +                      a   �  *         ����b   +  �         	   ����   O   �     
      ����P   a   �              ����                        ����                        ����                        ����                        ����                        ����            !                +      !               '  �            ����(  +  �  !      	   ����     �  !   
      ����  '  �              ����                        ����                        ����                        ����                        ����                        ����            (                +      *               >   �  (         ����?   +  �         	   ����      �     
            >   �              ����                        ����                        ����                        ����                     ����   1   �           ����2   >   �              ����                        ����                        ����                        ����                            +      *               �   �           �����   +  �        	   ����   �   �  2   
      �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �           �����   +  �              ����                        ����                        ����                        ����                            +      ,         ����      �                 +  �              ����                        ����            $      	         ^   �     
         _   +  �  %         ����      �  *               ^   �           ����_   �   �              �   +  �              ����                        ����                     �����   �   �           �����   +  �              ����                        ����            *         ����   2   �           ����3   ^   �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            $                +      $         ����   <   �  $         ����=   +  �              ����                        ����                        ����                        ����                             +                ����      �  '               +  �              ����                        ����                  	         T   �      
      ����U   +  �  $         ����   N   �  2         ����O   T   �              ����                        ����                        ����                        ����                        ����                        ����            -                +      -         ����   �   �  .         �����   +  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �        	   ����      �     
      ����   �   �              ����                        ����                        ����                        ����                        ����                        ����                            +               ����   �   �              �   +  �              ����                        ����                  	   �����   &  �      
      ����'  +  �              ����                        ����                        ����                        ����            !                +                     &  �            ����'  +    !      	   ����            
            &                ����                        ����                        ����                        ����                     ����        2         ����!  &                ����                        ����                        ����                        ����            *                +      -               p     *         ����q   +          	   ����   `     +   
      ����a   p                 ����                        ����                        ����                        ����                        ����                        ����                            +                     �   	           �����   +          	   ����   P   
  '   
         Q   �                 ����                        ����                        ����                        ����            /         ����Q   �     ,         �����   �                 ����                        ����                        ����                        ����                            +                      �              �����   +           	   ����            
      ����   �                 ����                        ����                        ����                        ����                        ����                        ����                            +      )         ����        *               +                ����                        ����            *      	   ����   p     !   
      ����q   +                ����                        ����                        ����                        ����            	                +      	         ����   
             ����  +                ����                        ����                        ����                        ����                            +               ����   j                 k   +                ����                        ����                  	   ����k          
           +                ����                        ����                      ����               ����  +                ����                        ����                        ����                        ����                            +                     �              �����   +  $        	         N      *   
      ����O   �   #              ����                        ����                     ����   )   !           ����*   N   "              ����                        ����                        ����                        ����                        ����                        ����            1                +               ����   �   %  1         �����   +  &              ����                        ����                        ����                        ����                            +               ����   t   '              u   +  (              ����                        ����            !      	      u   �   )     
      �����   +  ,           ����u   �   *  !         �����   �   +              ����                        ����                        ����                        ����                        ����                        ����                            +                     �   -           �����   +  0  "      	   ����   �   .     
      �����   �   /              ����                        ����                        ����                        ����                        ����                        ����                            +      +               �   1           �����   +  6  *      	         �   2      
      �����   �   5              ����                        ����            *         ����      3  *         ����    �   4              ����                        ����                        ����                        ����                        ����                        ����            '                +               ����     7  	              +  8              ����                        ����                  	   ����    9  	   
      ����   +  :              ����                        ����                        ����                        ����                            +      2         ����   p   ;              q   +  <              ����                        ����            !      	      q     =     
      ����  +  D              q   �   >           �����     C              ����                        ����            )            q   �   ?  !         �����   �   B              ����                        ����            )         ����q   �   @            �����   �   A              ����                        ����                        ����                        ����                        ����                        ����            ,                +      0               �   E  #         �����   +  H        	   ����   �   F  0   
      �����   �   G              ����                        ����                        ����                        ����                        ����                        ����            0                +                     '  I            ����(  +  R  0      	         o   J     
         p   '  M              ����                        ����            +         ����   g   K  0         ����h   o   L  2         ����p   u   N              v   '  O              ����                        ����            1         ����v   {   P           ����|   '  Q              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            (                +               ����   =   S              >   +  T              ����                        ����                  	   ����>   L   U     
      ����M   +  V              ����                        ����                        ����                        ����                            +      ,                  W           ����   +  Z         	   ����      X  ,   
      ����      Y              ����                        ����                        ����                        ����                        ����                        ����                            +                ����      [  0               +  \              ����                        ����                  	         $  ]  '   
      ����%  +  f  0         ����   !   ^  %            "   $  _              ����                        ����                        ����                        ����            0         	   "   D   `  %         	   E   $  c           ����"   ;   a           ����<   D   b  0         ����E   �   d  0         �����   $  e              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����            0                +                     %  g  2         ����&  +  j        	   ����   �   h     
      �����   %  i              ����                        ����                        ����                        ����                        ����                        ����                            *               ����   O   k              P   *  l              ����                        ����                  	   ����P     m     
           *  n              ����                        ����                     ����    o           ����  *  p              ����                        ����                        ����                        ����            *                +      *         ����   �   q  *         �����   +  r              ����                        ����                        ����                        ����                            *                     �   s           �����   *  ~  	      	         C   t     
         D   �   w              ����                        ����                      ����      u  	         ����   C   v              D   }   x              ~   �   {           ����D   w   y  2         ����x   }   z  1         ����~   �   |            �����   �   }              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            *               ����   
                    *  �              ����                        ����                  	   ����      �     
      ����  *  �              ����                        ����                        ����                        ����            $                +                ����      �           ����   +  �              ����                        ����                        ����                        ����                            +                       �                +  �        	           �      
      ����    �                '  �            ����(  +  �           ����   �   �           �����     �              ����                        ����            #         ����    �           ����  '  �              ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                        ����                            *      $         ����   �   �           �����   *  �              ����                        ����                        ����                        ����                            +                     �   �           �����   +  �  $      	         �   �     
      �����   �   �              ����                        ����            '         ����   �   �  $         �����   �   �              ����                        ����                        ����                        ����                        ����                        ����                                        ��m���?4'�'8S@WG��Љ@      �?�uT5A��?��DJ�@        �a�/�?      -@�l�� @        '<�ߠ��?�s�^o @����R�%@        Sc��|�?��C�lG@h/����.@        ��7�v��?p%;61@"""""@        ����o�?�;k�]h@s�H;V@        �VNx���?      '@j'p'p@        ��ݮ�?                        �"Qj�a�?                ��yVQQ@      S@                �TWέ�?      @                ��%|��?      @                ��[?"��      @                ��%|��?      @                ��[?"��      @                ?�;�S�      d@                ��e�U@      @                        �u�y��?      )@蘡X-�"@        �]+'<�?                ��ѡ%�      &@                ��a�+�&@      ;@                PE��w�      @                L��N��.@      7@⪲�`�?�N�B�[@              �?�ŊL�?Qb�(,@        }�(5�0�?�Ǻ��@l�fOS�@        ݮ���?     �<@���j(�&@        *.�u��?     @B@�+��n"@        )5�0ȧ?                )�SsH@     �S@                Dg̒8K@      K@      �?��^�
@        ��o���?      N@\s*�@        �|�(5��?                �v*���      @                (�3L{^$@      $@                l\;5�?      @                �^�֧&T�     �\@                ��ɣ.X�      @@                zV�V@      @.�o��%�?���PX@              �?��^�?�M���s@        �۵r�3�?     �=@�X�[�	@        �H�{��?L���|�?�ĝ�4%@        �0���?��鲘��?9B[�@        UUUUUU�?                0FFU@     @W@                 ���M?      @��W���?;�W�o�@        $J�=��?                        ;ڼOqɐ?U��7 �?�`p�b\@        �Y@�H��?j�t�M@IP�A�@        #Qj�a�?                ��p�m�S�     �d@                �sbD2�@      @                ��p�m�S�     �d@                �sbD2�@      @      *@                �Y@�H��?�y�t��?
e�?        �Y@�H��?                �!��\��      @                "Г'& @      @                �.���      @                +���
@��       @                T�C�e(@      @                V��X!@      @2��Y��?	c<��W@              �??�m��?���T-@        ��Y@�H�?��x�@ļɵ @        ��L�n�?     �W@v���=�#@        ��!XG�?˄_���?                #Qj�a�?�r.�5@��a�(�@        [9���?      )@s�v��@        F����,�?�"��J��?�+�[~@        e���}�?�҇.���?                XG��).�?                ���#�X�     �d@                X_�^���      *@                �.Q'Z�     �c@                �x���      *@                2�Q��Y�      e@                n����0�      @                (�".@      ;@                �a��׳�      &@                ��[��      @                ��[Y��N@      R@��d�z�?#�w�W@              �?Y���-�?�mi�b~@        I�{��?�%PV@W��r֠@        o��	���?                �k<RL�     �^@                xHV���     �K@                �.7$��2@     �A@                }�C�45S@     �U@H�}8g�?Z$��Y�V@              �?���|\��?�/Q�/0@        �ߠ۵r�?�@���
@��H�R@        Z@�H��?->�x�?��� � @        �n��	�?�bb�q@Ԡԏe-	@        ��L�n�?                Ga<�LD@     �Q@                ��%���D@     �G@                ծʭ�
G�     �X@                �;ؚ��C�      L@                HSO�0@      6@                �x\!e�@      @
ףp=��?
I�Z	8W@              �? �4��?�M@        �:ڼOq�?䥛� ��?j���Q@        ~�K�`�?                Q7�̈́�T�     @e@                :�HE�	@      @R�8��a�?�S�@        [9���?\*��{@��ڄ��?        '<�ߠ��?R���AD@�o�А@        ���:�?                        �"Qj�a�?                ��	�R@     �V@                ��,H���?      @                ���]¹�      @                ��s�(�*@      5@                ���]¹�      @                ��s�(�*@      5@�n����?d-R���[@              �?Ԛ��(�?�[�3!@        �{���?n��J���?"J&:�	%@        ��	��7�?                S�N�T�     �a@                >1l��      E@                �a�/�@      9@                �ߝ�:�T@     �V@��G�`�?�>�g]�W@              �?\ A�c��?�	�W$@        1��R�?       @D�`g��!@        ��o��Z�?t�3���?�t�@        f�"Q�?ꕲql�?�4c{��?        #Qj�a�?                        �k�g�{?���~�z�?�X��_@        �S\2��?                ?-��(�T�     @b@                �,�֩�      5@                �Vۡ@      @                �<� @      @                �Vۡ@      @                �<� @      @j���vD�?�}�M�@        )5�0ȧ?      #@M5e}��%@        J�=���?                        XG��).�?                        �"Qj�a�?     �0@��+	�@        XG��).�?      @��r1��?        _$J�=��?      @[��	o!�?        ;ڼOqɠ?��N�`]@;��ֽ{�?        ;ڼOqɐ?                4�#
� @      .@                ����*S@      T@                �O���?      @                
�:��j@      @                �NL�      @                .{=|g�      @                �NL�      @                .{=|g�      @                �NL�      @                .{=|g�      @���	���?v�Ʀ�R@              �?3P���?�X��(\@        &C��6��?������@HhnzcG@        �y��!�?      ?@�g�w�#$@        �E�����?�Y/�r��?�P��|@        ��|�(5�?                ��#�0@      B@                �[,�4P@     �T@                ��⫰tM�      ^@                ��Aǆ�@      @                �-��?      H@                �]HV��      @d���&�?�Sy�F;X@              �?�} R�8�?y=[�3s%@        I�{��?�_�5�@נ!�NG@        o��	���?                �0,��Q�     �_@                ��3�!��      M@                p��h��1@     �A@                ���N�Q@      T@d�����?u}�h�X@              �?r�t����?8����,@        ��o��Z�?�6�ُ@�u@        �, _$J�?     �=@�w�)� @        ��Rc�?'N�w(��?�P��ٌ@        �Y@�H��?t��m��?na�� @        �]+'<��?:X��0��?Ȇ�$Ao�?        �����?     �1@%��2@��_�s̿�ݮ��?                        ������?                n8�[�@      @                ��' ��?      @                \�E#��2�      H@                \p`�P�     �T@                \�E#��2�      H@                \p`�P�     �T@                �]�!*2%@     �J@                $c�Ж�8@      <@                B�%J�jL@     �O@                ���j�@       @�#�G[�?�Ywm��O@              �?;�O��.�?���jH�"@        �, _$J�?_�L�j@��>Ҹ@        x��A�k�?                �Ff,�R�      h@                �����@      @                �QI�t$@      B@                7��J@     @P@k��c�?˛�k�BX@              �? ���Y��?X-���,.@        �Y@�H��?\���(�<@4�]���!@        �L�n��?      @� ��%�@        �`mާ�? �rh�]A@C��NY�@        �/�Ʈ?                l�G-�Y�      @                &�5:V@     �^@                +V��J�?      *@                ��t_�V�     �a@                � .��      @                �o���%@      ,@~�:p�H�?�;iz)�T@              �?���g?R�?�qg�`�3@        �, _$J�?p=
ףPB@&-���@        x��A�k�?���מY�?��=�@        ��Y@�H�?�w��#��?�����?        #Qj�a�?                �dX�E�ҿ      @                �ӫ�xdT@     @Y@     �:@�(}��@        $J�=��?U0*���?��8��<@        j�a�/�?                �tfU�@      @                W�%�$�@      @                (��u�S�     �b@                �߫��b@      ,@                �_OK@      *@                9ݧ��      @^c��ޚ�?^�6��R@              �?+����?=�/�$<'@        ������?�A`��i@5�]�v�@        mާ�d�?      D@���[@        I�{��?��kCe@��>�/��?        �/�ƞ?                uΓ���R@     @Z@                !-�r]��      @     �A@�7ps��@        �n��	�?+����L@�#$� @        $J�=��?                �je��p@      @                [�<�?      @                N��IM�     �_@                �11�M,�      .@                /d��4!@      5@                �=�)v#�      3@���e%�?�W:Q@              �?�h㈵��?ؖm�2@        �۵r�3�?      @y���@        �H�{��?                �	�CK�T�     �e@                u�8��'&@      B@                �	T����      @                [W��g�O@      V@ZLl>���?����A�R@              �?N֨�h4�?)K0~�H@        �6�S\2�?jo��ɔ@�O��@        �!XG��?      @�,[��@        UUUUUU�?T �g���?ς��S�@        ��Rc�?                ,7��� @      8@                �'��
(S@      X@                        �"Qj�a�?     �1@*-����@        &C��6��?                iK��@      ,@                �����3�     �S@                iK��@      ,@                �����3�     �S@                �u��/2�      4@                w�s��?:�      O@B	3m�
�?���I�Q@              �?P�2�ˢ�?�矊7@        ~�K�`�?��#bJd�?�6�n�9@        �h�>��?     �;@m/[p�@        �k�g��?+~����?I3��p%�?        j�a�/�?                ���!�;@     �I@                �?�[��D@     �G@                й�+��N�      Z@                ���ob/�      U@                �[Te>@      @                |Ӌx�@      @I.�!���?�5���P@              �?g��j+��?����(@        �a�/�?     �N@��މ@        '<�ߠ��?G�ŧ ��?;���+@        �k�g��?kH�c��?��O� h�?        Sc��|�?     �A@JO$�Fc@        ������?                        �k�g��?7�ُ��?����b�@        �������?^�c@�z�?S{	���?        ������?                �ȟ���?      @                .U`�q�@      @     �=@~8r@        ��!XG�?F����E@��bn�@        v�y���?                [�V���?      $@                $�"�>KO@      U@                        ;ڼOqɐ?�������?                �u�y��?                        �"Qj�a�?k}�Жs�?іr�s�?        F����,�?                wc���      @                n���P@     �S@                �̸c�� @      0@                �k/$�K@     �O@                �̸c�� @      0@                �k/$�K@     �O@                ���f�<@      @@                �&\�A@     �G@      )@�:�_�A@        f�"Q�?                        �"Qj�a�?                �z�(��      @                �<��p!�      "@                ��'n{�C�     �K@                �|�FG�@�     �]@                ��'n{�C�     �K@                �|�FG�@�     �]@�x�S�?��Q��FS@              �?     �Y@5^�E��$@        e���}�?������1@{�1�-&@        7�S\2�?                �/X4��S�     �c@                bO,�<�@      2@                ѐ#�k�      @                ��pv�S@     �]@^�,σ��?�S�k�R@              �?      @�4��� (@        ~�K�`�?m����">@KN�?]�%@        �h�>��?      6@ټ�F·@        j�a�/�?�B�O���?WL��M�@        �k�g��?                        ��ݮ��?K<�l�U@'i�`fd�?        ��|�(�?                (.Ŀ��?      @                �нs+�@      @�m�2�?��~���@        ڼOq��?     @@@B5�[�@        )5�0��?                %p�bg�L�     �_@                6�����      K@                ���̝�S@     @W@                �|W���@      &@     �8@m�[H�@        Z@�H��?                        �/�Ǝ?      T@�z���(,@        ����o�?      ,@m���@@        �}�K�`�?�N�z1T�?�~h@        ��E�Ը?}iƢ�?                #Qj�a�?����Qr�?�tI
��@        �k�g��?��H����?�J>:�V�?        �/�ƞ?                �Q����?      @                Gr.���3�      9@                �m��)�      6@                ��Q�N�      @                d�����      @                /��`'�?      @                ��<���	@      @                �LƄ�@      @                d�����.�      N@                ����3�F�      O@                d�����.�      N@                ����3�F�      O@��^�?�.i�'0R@              �?N�St$�?���,b0@        �0���?��HP�?�`�]@        ��o���?                1���GVR�     `b@                r\>n��      =@V�F摿�?���R	@        �Y@�H��?Á�,`�?�n0i�@        ��Y@�H�?������?cQ����?        �k�g��?��b('�?����4�$@        ��ݮ��?=
ףp�N@��m�K@        UUUUUU�?ƿϸp�@��P��?        �d����?      2@�*���@        ��ݮ��?T㥛�|Z@`)�'�:�?        �����?                D��2*K@     �O@                �AP��c�?      @                        ��ݮ��?                        ��ݮ��?                ���l'#@      &@                ވ��4�?      @                ���l'#@      &@                ވ��4�?      @                ���l'#@      &@                ވ��4�?      @                ����@      @                �_�����?      @     �9@s?��>�@        �}�K�`�?     �4@Տ����j?        ��ݮ��?:3P?�?��8��?        �/�ƞ?      *@                �k�g��?                �{vg�?@      @                GM/V,�@      @                M���R��      @                �íb�l�      @                ;=�u@ �      @                ͈�y8B�      @k��c�?���%�S@              �?�(�~�?�3I3�Q$@        �Y@�H��?�|?5^��?��gQ�@        �L�n��?     �Z@l����5"@        ���:�?                        �"Qj�a�?                ;+G5�@      ?@                ���t�&S@     @Z@     �:@S���@        ��D��?�4S�?                j�a�/�?                aX>��R�      c@                Z���&(@      @     �8@K'id�@        �/�Ʈ?     �R@��un@,ւ���.�u�y�?                �?��R�      b@                eC�:���      @                �GD��@      $@                *} �y0�      @                �; ��xS�     @`@                D	�m�+�?      @@�Ŋ��?0D3��N@              �?     �D@��NyX'@        �������?����@b��@        �������?c�tv2x�?&"��p�&@        F����,�?     @G@�r�Z�@        &C��6�?                ]�!L��P@      Z@                �v|����      @                ! & �R�     �d@                )�>��t@      @                ��|td�@      @                �$q�B��?      (@V�`��?��z�O�R@              �?RI��&��?"����@        ~�K�`�?|�w�@�	x����?        �h�>��?      V@;�9u� @        ܵr�3��?��s�/�?�	@�U�@        @�H�{�?                >�s �R@     @X@                .� a�V�?      @      �?�:l��@        ��7�v��?^����?                ������?333333F@��°� @        �"Qj�a�?                        ;ڼOqɐ?                n��Vme�?      @                `SK�<�O�     �`@                S���K�      `@                 �Sb��      @                �rC�}�!�      ,@                �Ņ��"@      C@                �rC�}�!�      ,@                �Ņ��"@      C@�|?5^��?�ݲ1��P@              �?9�ߡ(��?�����@        ܵr�3��?�����@)���:�?        I�{��?      �?�L���m@        ���Y@��?333333F@���%=�!@        ������?                �����0@      B@                �1-�@I@      Q@                        ��ݮ��?      -@/?r�@        �y��!�?�p=
׳C@R���?        �"Qj�a�?%��CkI@Ed��@        �/�ƾ?                2{�;� �      "@                 EAH�8��      @                _�Y�@      @                ��_d���?      9@                _�Y�@      @                ��_d���?      9@                �l-�,�?      ,@                -�E�vQ�     �`@䥛� ��?��q���E@              �?��I�r�?���2��)@        �a�/�?,e�X�@��B$���?        '<�ߠ��?      -@!6��Z#@        �6�S\2�?w��N#��?Q����?        �k�g��?                vE��H@      S@                 ���D��?      @��bb� @̎N\�`"@        ��D��?2r���?�,���@        �g�t��?                "GF	�@      @                ]L��ͪ@      @                Ʀ���L�     �V@                �`��o@       @                �I
��1�     @U@                �醵�@      5@ZLl>���?\)�/@�J@              �?8�����?�y�QH@        �6�S\2�?�%PV@�WY�� @        �!XG��?R'�����?�9��v@        �E����?T �g���?,�z��@        {���?                �aJ*@     �@@                2:Y��DJ@     �R@                &}��]G�      U@                ��\��@      "@                P����@      5@                o&oo�0�     @S@S�
c��?V�!��Q@              �?      @�>�o[#@        �������?b֋����?��A�)�@        �������?      &@-�Oa@        �Y@�H��?     �8@�QB7G@        ާ�d��?                �Pw���@      <@                �חw�
Q@      Z@                g�~"H��      @                ����x�@      @                �Dr|&�L�      U@                E�P��}2�     �Q@���{��?��M8��I@              �?d�]K�G�?dP!@        �u�y���?     �4@7]I�S�@        ���:�?�S:X�g�?P!2%�@        *.�u��?      *@~���	@        �u�y��?                @��ۙk@      @@                ���Q�O@      V@                ��)�I�     `d@                !��J%�      @                �Fܚ���      @                š��2�@      @�|?5^��?�ql�7J@              �?�]P�r�?���q��*@        ܵr�3��?��ʡEL@�X�M�@        I�{��?     �X@�m��Iq@        ��Y@�H�?�T�t<f�?�o=^���?        ��!XG�?��"�-@%�9t�@        �����?�C�l��h@�P#4@        �f�"�?      9@�p!I1@        $J�=��?      _@<���FP	@        j�a�/�?                �[�"@      ,@                ��r��߿      @     �1@~�����@�#�k<������o�?     �?@�K[/�'�?        XG��).�?                
ŢF@      ,@                �e����       @      $@0��)��@        WNx��A�?      @�o�u`@        2�h�>�?                XO��d@      &@                J%QX���      @                ��e��      @                C����?      @                ��H�K@     �S@                ����b�?      @      6@�I	Ӌ�?        ��ݮ�?     �7@��@�@        ާ�d��?                        XG��).�?����~$�?�����?X��	6ٿ�).�u�?                D�z��|@      @                ���@Q�     �W@                c�%���F�     @Q@                �^T#��7�      :@                R�=�|���      @                ��V��A!�      $@      D@����@        Sc��|�?     @C@�I�d�� @        j�a�/�?                7�͆k�"�      *@                �8rtz��      "@      )@!LC�@        �k�g��?                        ;ڼOqɐ?                [�_�*�      @                ��R�lI$@      &@                [�_�*�      @                ��R�lI$@      &@=,Ԛ���?�f��M@              �?�=���d�?��R{@$@        ������?��&SE�?��U��@        mާ�d�?�D����?�3�_Z<@        l�g��?��:���?                �k�g��?��	��C@Q�VԘ@        XG��).�?.9(a�!@�8S��{�?        .�u�y�?                D��"\K�      f@                ��OV�'�      ,@                � B3�P�      f@                 q3u�m�?      *@                ��5j@      7@                �Էs2@      @                3�����J@     @Q@                ���U�u�?      @2��PN��?dj׵'2P@              �?PjM��?�r����-@        I�{��?Hm��~��?zp����@        o��	���?     @@@K��.�q@        i�>�%C�?��x�@�W�e�@        �ݮ��?                e42
(@      A@                g��`�K@     �R@     �;@��l٘	@        >��E��?      Q@�X�Hk@J�j�u���)5�0��?                uW^�ݟ	@      ?@                �3J��@      @                �-��6~;�     �P@                q�h!��?      4@                ����_�G�     �O@                �kTL���?      @W�c#��?����N@              �?     �<@�����^&@        ��|�(�?��x�@w����?        ��ݮ�?                �/��[P�     �e@                ͳ�^b� @      8@                �>�a�%@      8@                AD�-)�L@     @S@���=�$�?�����H@              �?     @H@�����%@        ��|�(5�?     �I@T�(�@        ��ݮ��?�Cn���?+����#@        �n��	��?     �J@*0_�@        �"Qj�a�?�<,Ԛ��?                ������?�(\��yc@��a{�?        �=��E�?�-�l�I�?>����c
@�(^gE����ݮ��?      %@��N��@        ��ݮ��?                �aF|��@      @                N��~D�@      &@                �	l��J�     @e@                ���E��%�      *@                5�p���      @                ��^�g� @      $@                ��s�+H
@      @                ^G��@      "@                a���L@      R@                �dl��@      "@� �> i�?�%���C@              �? ����}�?���*=� @        }�(5�0�?1��*d�?�p�N��&@        ݮ���?                ����NG�     �c@                �x* ��@      1@     @@@;e�}i '@        ���Y@��?                        �k�g��?                ¨��n�Q@     �]@                k�a?F��      @                ¨��n�Q@     �]@                k�a?F��      @��n��?��WN�EL@              �?�� ���?{����o$@        ��|�(5�?��n @����\@        ��ݮ��?\Υ��L @̥:؞�@        �H�{��?�E|'f��?                ��ݮ��?     �6@�����@        ��f��?                        ��ݮ��?��N�`}�?��YJ�@        �۵r��?Mu�T�?~S%>�?        �}�K�`�?                rh��P�     �e@                \2L��@      "@f�c]��?Pmi� "@        e���}�?�K�����?��>5�?        ��Y@�H�?                ���?      @                3�m��/@      @�£��@^B�m,m@        �/�ƞ?      O@a�wk�?        �����?                �N/By��?      $@                ���pQ@      X@                ���2_�      @                x��Z��@      @                ���PVN@     �S@                ʢ��{�@      1@      @v���@        {��D�?������?�a=����?        ��ݮ��?                ������      @                �'%�;��      @                �V[��@      @                �b-#Q�     �b@                n�aZ�@      @                ���|-��?      @�x�S�?�9x"zI@              �?     �Y@M��@��*@        e���}�?��ek��?�gd]d�@        7�S\2�?                �o�%�O�     `c@                z�U5�!@      .@                wtI6��@      @@                �rb[I�N@     @X@���+�?#�f+�E@              �?�+H3��?$�@ߘk@        I�{��?!Y�n�@*�0̥��?        o��	���?��(\��?@t�C��!@        ��:��?0��{���?���Pҵ@        �"Qj�a�?                A-�/@      D@                ��>vJ@     �T@      E@��X�)@        )5�0ȷ?��Q���?�$����?        �	��7��?"���?�r0D�"�?        �����?z�Cn�[�?-���N#@        �7�v���?��:�?                �u�y��?/�$�7@�V�r��?        ��7�v��?                ���lA�      W@                ��� )�'�      0@                )KϨ�F�     �Y@                �eIubs�      @                \b����?      @                �Q$"@       @                �z�N@      @                �D��@      @                �D�W�s�      *@                \o�5@      ?@����F�?�4Y]�WB@              �?��x�&1�?�g7mcH&@        B�k�g�?v��y���?6��_�@        }�(5�0�?                l���M�      e@                �z���@      @                �!+�F�@      D@                �Vm_�F@      U@d]�F��?�M�>kbI@              �?d�w��?!�C�'@        <�ߠ۵�?K�h��?�4uݭR&@        �Y@�H��?     �D@)��N@        [9���?�;k�]��?��&��@        ;ڼOq��?                ���ᛵ�?     �D@                �h~�J@      T@                �3э&Q�     �[@                ��/W��      <@                a���Ē#@      7@                o#E7�      1@V�`��?�����G@              �?Է�鲘�?W��C��#@        ~�K�`�?(�$�I@'��/_a�?        �h�>��?     �Y@0��m$�@        �Rc���?���:�?                ��ݮ��?                �_0��0@      E@                2�m�xGD@      N@     �<@�л�l@        �0���?      9@��TX�% @        .�u�y�?                Y̸S�N�      g@                lz+��?      @                �&~���K�     �Y@                =����U%�     �P@                        ������?      0@Y�d�\m@        ������?                ��U���      @                9e�qi#@      0@      /@                XG��).�?/�Xniu�?�"a(k٫?        �}�K�`�?                ��Cs˨@      @                ��pW)@      &@                #%|�|@      @                
��X�@      @��҇.h�?����@F@              �?     �9@��M¨�
@        ��|�(5�? o�ŏ�?v��Qu&@        ��A�k��?                �K-���<�      C@                �jN�dc1�      H@J��Z���?��^��@        j�a�/�?R���AD@5�{*M)@        �!XG��?                ؖ�W
�#@      ,@                ���賁�     �R@                ���۰^�      (@                �Y��g3Q@      \@F���j�?� ��B@              �?���+�?<o��g?+@        �=��E�?      <@&E=`�'@        �g�t�?�����l3@�˓��7$@        ���Y@��?     �:@4���?@        @�H�{�?      @j �B�e$@        M�n���?     @@@�/��M�?        �Y@�H��?                s]Ҍ��@      @                ��7��P�      c@                p�[=�O�      @                ��R&#@      $@                �&�����      @                ����N@     �]@                �� G;���      @                ��&2G%�      @"�uq��?��{#ȵG@              �?^�}t� @Y��Q�@        s�3���?�G�z$H@=�ew`@        {���?                G載�NP�     `h@                �K�6=@      &@                B�����      "@                ��6%9K@      U@~�:p�H�?xE�P%4J@              �?l}�Ж��?�KY5&@        �, _$J�?     �W@��y��@        x��A�k�?                ���MP�P�     @g@                �^~j8�@      @                �����aN@     @Y@                �Og�����      @_F�����?��,�.>@              �?���N��?�_C�!%@        {���?F*�-9�?~�^d�I�?        �	��7��?                ��j��QE�      g@                xO��p!@      &@                �5�I�@       @                �R�&�E@     �W@���e%�?	 �8�F@              �?      @gqy%�"@        �۵r�3�?     �P@'z;�aV@        �H�{��?       @��yO���?        �"Qj�a�?     @A@UUA!�"@        �Rc���?                �[��3�J@     @W@                ���1VK@      6@                @D�wr��?      @                �'�	��@      @8��d���?%� �Y@         _$J�=�?                        ;ڼOqɀ?                lLBD�!Q�     �d@                ���&s@      @                lLBD�!Q�     �d@                ���&s@      @"��u���?��-1&H@              �?     �Y@p	l�*@        ������?��uz@<��D&�@        mާ�d�?�=���d�?��NZ�%@        ��o���?      ]@sN���@        ����o�?                %wR!t�M@     �W@                ���      @                �(!�NR�      e@                :��E�@      "@                :H���v@       @                �Pꊨ�@      .@��~��L�?����E@              �?^.�;1k�?�y�M�@        B�k�g�?      @�u`�@        }�(5�0�?                Z��*W8�     �Y@                P��7hGA�     �Q@                        )5�0ȗ?�n��\g�?���j/@        *.�u��?                �&
T�      @                Pd�:yM@     �^@�*5{�U�?o&cq�@        ��E���?                        �k�g��?��A�&�?�0��Y	@        �����?\���(�E@M����?        �Y@�H��?                l��ɎC0@     �J@                /�	XF@     @P@                ������0@      A@                 �G�y�ؿ      3@                 h�O�Q�?      @                7�r�e5F@      O@2���#�?pu�W`g@@              �?     �X@'(�YI#@        C��6�S�?�@+0d�@#V4�#�@        z��!X�?                ��_uTL�      g@                ۸/#�@      @                b�4 Gy#@     �H@                BJ'B@      N@�������?קa��-H@              �?�����?����С(@        J�=���?      5@2��ﳔ@        l�g��?                H�D��N�      h@                Q�>�@      "@                Ļ�.��?       @                ���`{�L@     �V@n��S�?�w���E@              �?     �8@�[\h8 @        C��6�S�?��x�@� �U�@        z��!X�?                O�z�_oN�     �b@                I>��g@     �E@                ��{C��@      >@                �@k{�G@     @S@��m���?.��&D@              �?     �Y@p��a�.'@        �a�/�?L7�A`�;@#"��T@        '<�ߠ��?                g}m�"L�     �d@                a6jQ�#@      9@                �\����      @                ��P��L@      Z@��4)��?t}ʺeQA@              �?l�`q8��?��Q��$@        ���}�K�?33333�h@b�Q��@        T\2�h�?�'��?M��RI@        �]+'<�?\w�T���?�b{��3@        @�H�{�?                �Se{ֱJ@     �V@                �t���      @                ����C�      d@                X�w "�      $@                �Į�����      2@                Ƙ�*��(@      .@
pU��?䁣��@@              �?�F�?�?��ۯq�@        �S\2��?     �=@g�˘4"@        "XG��)�?                �P�]9�     @\@                ��z��G9�     �I@       @�ŔV��@        ��:��?�
p�@�"�K��@        ������?                        �k�g�{?�5���@���W��@~I�ȩ}?f�"Qj�?                ��s�t��      @                :4"�?�?      @                ��s�t��      @                :4"�?�?      @                pE��N@     @]@                �%��*�      @R�i>"�?��m�D@              �?     �K@�1'�Ĺ%@        �۵r�3�?�je�/@Չ:|q�?        �H�{��?     @A@�/��J|@        {���?�B�O���?                ������?                c��9@     �N@                !awK�8@     �B@                �[�RgM�     `b@                �,���      H@                q��P�     �f@                ��^�i@      *@X��0_��?�%�QQ"D@              �?     �8@�+�|�!@        [9���?F����E@f��t(�@        J�=���?     @^@ڸ�׾�@        ��Rc�?!Y�n�?���	�G	@        .�u�y�?                ew Ӵ�?      $@                �$Η MJ@     @W@      J@���@�@d��U���B�k�g�?                        ������?                ��Ik�"@      .@                �>#����      @     �D@�`��n@        �f�"�?�V`���?V$�dG�?        ��Y@�H�?                8�D��&J�     @d@                ��M���$�      &@                �By��eL�      a@                U����@      :@                ��[�<�      @                �=��~<�      @�������?��V�@@              �?      @߳y"5,@        J�=���?�9]K@ƥ�&H @        l�g��?     �2@��P��>�?        j�a�/�?     �6@���1.@        �n��	��?                i{0�A�H@     @U@                 ��Hs��      @                3��֥@      @                �f�j޷@      @                �@#�K�B�     �V@                ޾��+� �     �[@�1��o�?.Wȴ\A@              �?v�k�F=�?Ad�V��@        ��f�?_�L�j@��cP@        ܵr�3��?                �3��nC�     �^@                B�_QG�     �C@l	��gs�??��e�_@        ��:��?)\���x[@�����	@        ����, �?                �感�� @      *@                ����t%@     �L@�) �3��?&
��B��?        q�����?                        �Y@�H��?                5f�@      @                �4���B@      M@                5f�@      @                �4���B@      M@.�o��%�?a���P"G@              �?      @�1澫%@        �۵r�3�?��+e�@9x8���
@        �H�{��?     �B@#GM��X@        #Qj�a�?     �7@��%�|�@        �6�S\2�?                �m��rN@      [@                x0�!a��      @     �:@�嶺cM�?        �"Qj�a�?                        ��ݮ��?      /@}�!�4\@        ��f��?.�l�IF�?�C(��0@        x��A�k�?                ��v秚@      @                �FC�FY@      @                ��v秚@      @                �FC�FY@      @                ���<%�&�      C@                �j��ϰ<�      E@     �:@����@        �7�v���?     @@@��;�@        �]+'<�?     �6@��{"�y@        ��ݮ��?'�o|��?�h��@        C��6�S�?                M�͍s �      @                V�y�i
@      ,@                        ������?      /@                j�a�/�?     �@@�����o�?        �D����? �U+��?��d�  @        �"Qj�a�?                �3�611�      9@                 ��_+�     �@@                /m�jX�@      @                ���!��?      @                /m�jX�@      @                ���!��?      @                � P`kM	@      @                �?;E��?      @��s���?���ȕ�A@              �?     @O@a�l��?"@        �"Qj�a�?.�l�IF�?�ʡł@        �]+'<�?      9@@��!y� @32�uũ�����:�?     �:@! �~}S@        �7�v���?                >��)���      $@                ��MN3�E@     @T@                �V�G��Q�     �c@                k�g8 @      *@                ��)��      3@                �����&@      4@���e%�?c���	�A@              �?6Y����?���&�@        �۵r�3�?��+e�@' ��}@        �H�{��?*Ral!��?�
nr"�	@        ��7�v��?                        ;ڼOqɐ?                f�G2�I@     �Y@                ��P<�       @�Y��?�?}�,�ړ@        }�(5�0�?t$���� @��@        )5�0ȧ?                ;�$]E�      e@                ����&�      .@      @�W6P�@        ���:�?��kC��?97RE��?        �/�ƞ?                �[����%�      &@                �w��eӿ      @                �2�s�@      5@                ��R`J�     �a@                z{���-@      @                {?k����?      @V���n/�?9���Xi;@              �?�W�L���?>¶��,@        E���Y@�?��JvlD@��o��=�?        w���L�?      �?��\JɁ$@        ������?��k�U�?��5>�?        �Y@�H��?                G�
�V�6@     �N@                6n����3@      ?@                �+�AO�@       @                 �\�LM�     �f@                ��'�s%@      *@                �Oi����?      @��`�?�Ov�-:@              �?     �8@N���W#@        - _$J��?ףp=
Wa@�o�h�U@        ��A�k��?     �@@^q����!@        ��ݮ��?t�3�N�?����7@        .�u�y�?     @J@�a[.�@        #Qj�a�?�(\���@���4/�@        �]+'<�?��~�T$�?�"�ne�@        ^+'<���?     �3@�򊰃
@        ��ݮ�?                �1�����?      $@                �Q�ʙ@       @                �F�+F�     @c@                )�Y�"�      @                ��-�V@      9@                !���t1@      @                ���.6�E@     @Q@                ����#޿      @                I��z���      @                ��W�ў@      ,@I.�!���?��+&�@@              �?     �Y@����a�0@        �a�/�?      %@d"�7i@        '<�ߠ��?^�`7l�?�{0�0*@        7�S\2�?     �0@�����5@        ����o�?                .�*O�@      =@                ;�5�F@      S@��, �?gu(�J@              �?      2@��`��@        �y��!�?                4bi�.�      @                ��Q�P�*@      (@     �U@Ga�h�?D(�
��ݮ��?�����?                �/�ƞ?                �|�=��&@      ,@                ��E F��      @                �bs�z>M�     `a@                i�BA͌#�      (@                6�bq�CQ�     @b@                -DO����?      @�uT5A��?�i ��DA@              �?�Zd;�:@�i�ߐ�@        Sc��|�?���+�@��˾!^@        [9���?     @G@�ɵ�@        �Y@�H��?��(\��C@��Q��@        t�VNx��?                ��5���H@     �^@                yMI4����      @                n�9Y# @      .@                �n�S��      @                ��1�b�4�     �@@                �A#�Y�B�     @^@k��#�??A�h�tA@              �?     �=@ܗ8I��@        ��Rc�?
ףp=zF@�Xd�32@        �t�VN�?                �G`j�kL�     �a@                ri�ʇ@      @                �̒���%�      @@                Ǐ�/N@     �]@�=�$@��?�$��=@              �?     �5@�V3yp#"@        s�3���?     �;@��ש��@        {���?      �?����@        �t�VN�?     @X@��L�@        �h�>�%�?     �e@�P�f>�@        w���L�?                        ;ڼOqɐ?                P��:�?      @                ��*���E�     �Y@                &қ3r�@     �V@                @��p4�      @                /yF�̘I@     �V@                b5�)�:�      @                /yF�̘I@     �V@                b5�)�:�      @ܢ��$�?���Q�;@              �?�4�O��?�� %��@        Sc��|�?XV�����?� b	��@        [9���?                �/q)�7�     �_@                Ӕ��K4�     �B@                ���M@     �K@                �^@Y�vD@      T@DԷ�)�?��W$-=@              �?     �6@�c$�$@        t�VNx�?�z�G�F@�	jv��@        ��Rc�?      @����$@        �h�>��?      M@� 9:�@        4��]+�?x����,�?�����"@        ��Y@�H�?\���(�L@�%����?        ��}�K��?      -@�.�`D�@        @�H�{�?��:��?;a�%S!@        <�ߠ۵�?��$�?�i�&#@        mާ�d�?                        j�a�/�?��x��?ǖ*0���?        �Y@�H��?�X��@�?                �k�g��?                kvt��0#@      4@                .���B@      M@                ��I�U�@      @                �x�1@      @                �	��fP@      @                nؠ��@      @                        �Y@�H��?                        �"Qj�a�?      )@��2�� @        Sc��|�?5�8EGr�?                ��ݮ��?      !@�.�oD^@        �K�`m�?ףp=
�W@�A#�@        �۵r��?                yW�~D�     �R@                �����      @                yW�~D�     �R@                �����      @                yW�~D�     �R@                �����      @      -@�j�u��"@        *.�u��?      >@��=�Ę$@        ��6�S\�?                y�����(�      N@                T�3��H3@      I@?W[��l�?g4���?        �y��!�?     �2@�1�@        ��!XG�?     �B@��xE @        ;ڼOqɠ?      @5���@        C��6�S�?                �}_���      @                �0Ri�̿      @                        �k�g��?     �B@���6��?�!ur}��?��E�Ը?                ���)�      2@                (��>%	�      @     �1@�w�5�G@        &C��6�?     �@@U웎�@?        �}�K�`�?                w{���"@      >@                �N��N�       @                ��5�M6@      9@                R���'@      &@     �0@���4q@        ����o�?                        �k�g��?                <p�      @                и����      @      +@�ɑ��?        j�a�/�?��S��@@m�m�d@        )5�0ȧ?                MM��'@      @                @ݳ@帿      3@                %��~@      @                ��8��?      @                        XG��).�?      +@�E4����?        Sc��|�?                r�%7��@      @                �5�9R1�      ,@                �1A��}�      @                ���e+�?       @      )@gR$����?        ��!XG�?      9@K�9�7�@        ;ڼOqɰ?                �?���?�     �C@                V���[�?      @                PS�k�#�      (@                ������ �      @ףp=
E@��!�@        �Y@�H��?      F@�t�D̒�?        ��Y@�H�?                ��l����      @                %�r�@      @                 /y��      @                ?�R��	�      @Լ�I�?�zѧ(;@              �?8��m4@�?�!��?&@        �, _$J�?-���w?@������@        x��A�k�?     @K@�1�nYO@        ���, _�?���3KB�?ەv����?        �}�K�`�?                
?R���      @                `P�/�CF@      W@                ����bL�     �g@                #��u��@      "@                �{��z�@      @                d�^@      @���+�?D��g?@              �?�ѩ+��?��(:��@        I�{��?fk}���@�O���@        o��	���?                �W1�=HB�     �V@                ����~�.�      X@                ����	2@     �P@                �����9@      G@�P�fo @s�*�E�9@              �?�4c�tv�?�L4�#@        4��]+�?     �P@��\�@        ��D��?      @C<�@� @        UUUUUU�?�ŏ1��?i~ǣ2j�?        �}�K�`�?                ��V��LE@      S@                >MS��C�      (@                        )5�0ȗ?     @E@+��`@�8}`�ӿ������?                �-���@      @                >G���@      &@                �-���@      @                >G���@      &@                ���$_<L�      f@                z1��@      .@���խ~ @`�� a�9@              �?     �A@����Z�!@        WNx��A�?�e�--�?�Һ�
�@        Sc��|�?-`����?�@�x@'�p\Њȿ0��f�?     �9@:߲@�W@        ��L�n�?                C�g��?      *@                ��K/�vE@     �R@                �@�l�E�      a@                ��kʱ]�?      3@      (@٭��v$@        l�g��?     �;@�O[��A?        �Y@�H��?                �^6�φ/@      5@                `t�7>��      <@                㒜�u� �      @                �g)a
(�      @^�,σ��?�{tM,>@              �?\�C����?<c�ju�@        ~�K�`�?,e�X�@�>tdC�@        �h�>��?�7��d��?m앏�@        *.�u��?��מY�?٘#x��@        ��!XG�?                κ�A�C@      U@                ��<�6�      @                t��B�     �a@                �(��j�2�     �A@     �0@ʜ���@        �ݮ��?�Fw;S�?�G��Q@        @�H�{�?                        XG��).�?      7@|������?        )5�0ȧ?2 {����?9���@        j�a�/�?                        XG��).�?                ����      .@                ��/,���      @                ��_�[�?      @                ���be@      @                U����      $@                ����@      @                U����      $@                ����@      @��=�$ �?�2���:@              �?�HV1�?а��%}@        {��D�?     �=@"k���@        
��7�v�?N֨�h4�?�σ��@        �7�v���?                        ������?                4��p��I@      a@                �6DD�m�      @                #�>53�     �W@                %��h��:�     �L@                #�>53�     �W@                %��h��:�     �L@���e%�?�o:��@@              �?�ǘ���?�h�f"@        �۵r�3�?�z�G�F@�K3�	@        �H�{��?���m��?�o�6�@        �=��E�?     �0@����w� @        ��L�n�?                P����?      0@                <��j2�F@     �U@.�l�IF�?&�/[��@        �S\2��?��ʡE��?��{oi��?        ��ݮ�?��1ZG�?^M�LU�?        @�H�{�?     �B@���[I@        �"Qj�a�?                ����=@      @                ���A`@      &@     �2@���ə?        XG��).�?                        ��ݮ��?                �b�	�      @                e狩��      @                �b�	�      @                e狩��      @                �ɵ*[�I�     `a@                ����m�@      0@                {�����#�      $@                K��\c��      @�.n���?����@@              �? ��&N�@Yi�:��!@        ������?     �4@CT@!;x@        mާ�d�?��7��?<S�S�@        ڼOq��?{��㽪@.�k)?�?        �}�K�`�?                �e�s��?      1@                ��N�I@     �W@�4c�tv�?*X"&�q@        T\2�h�?�@H0��?�Q:,w�?        ������?                `��@      @                ��JU@      @                �4���;�      T@                ��
ۺ!�     @V@                @���tZ�      @                ��Zi-�      @��	my�?Ʒ�m�@@              �?�i>"��?�.�v@        ���}�K�?XV����@ba��3#	@        T\2�h�?                �����F�     �`@                ^j��$��     �Q@      /@��1���@        �=��E�?                        j�a�/�?                !�vx�?      .@                bSQ��E@     �S@                !�vx�?      .@                bSQ��E@     �S@��67�g�?��G��8@              �?     �V@y؟�O+@        �Z9���?����so�?Q=�e��?        $J�=��?      +@�ڱ@(@        �{���?\���(�H@�/���@        ��E�Ը?                	_R=*@     �D@                .����]:@      H@                �.�7+N�     �e@                ��ƪ� @      (@                �<�z?��      @                �8^ �x,@      1@K��>�?Ɠ&�2�<@              �?     �R@��P=q7#@        f�"Q�?      ?@ƌCG�#@        �3��]�?      6@=q���|	@        Sc��|�?      #@��$Ho�@        �Y@�H��?pB!a�?�?M��#�?        �����?                        ��ݮ��?                ��ȴS)@      G@                S�R�2B@     �R@                ��ȴS)@      G@                S�R�2B@     �R@                ���2��?      *@                �%��)�L�     �b@                �;�_03 @      @                �v�č�      @HĔH���?�~��N�7@              �?^F���j@��%I &@        ���o��?      @-���
@        ���, _�?� �t�?u ���r@        {���?V�F�?�?�'�>���?        ��Y@�H�?                �
�"���      @                Iřv�$E@     �S@      %@�W���@        �/���?�L��[@-�㗪@        ��f��?                ������@      @                �}2G �@      &@                �z�4�y@      @                ,�b���C�     �Y@                s�&�@      U@                q�����      $@����M"�?��6�7@              �?     @^@��_���#@        ��:��?^�D�
�?�@-)���?        ���}�K�?+���7�?H���ɻ @        ��]+'�?      R@�at���?        �"Qj�a�?                � ��Q|@      @                �Vq̰>@     �W@     �B@0[��8@��&��ȿ�3��]�?Z�����?                XG��).�?                �J�0
@      @                �;��@      @                Rq�:y:O�      b@                DDq!tٿ      E@                o �x��M�     �f@                H��P���      @���">�?�#d�cB@              �?      /@"��O|b@        Nx��A��?kH�c��?�
���o@        c��|��?                �����     �T@                �����E�     @X@                /�h���
�      "@                ��V���K@     �[@���Y@��_� 6@              �?�|~!�?	��'�f@        F����,�?      @�)t�_�?        �v���L�?Y��9��?y/����?        e���}�?jM��?��u�@        '<�ߠ��?                        ������?      @�b����?        ��7�v��?�je�/u�?�mǮ��?        XG��).�?�x�@e��?�Y�9�rx?        ������?T㥛Ġ�?�-�"ئ@        �۵r��?      -@U�B�"@        o��	���?     �Z@Q�|�D @        �]+'<ӿ?�m�2��? 7���h�?        �/�ƞ?      )@I� ����?        �Y@�H��?     �A@�xw�#@        �:ڼO�?                ��f}<@       @                7��hq�?      @�y�CnF�?,�I�!�@        ��ݮ�?     �0@6�[�f@        p��Z9�?���J�?���=^@        ��ݮ��?u��&�?�)ͬrq�?        )5�0ȧ?                        ;ڼOqɀ?��a����?<�ӊ��?        ��ݮ�?                _M�=���      @                9�e�W@      "@                ����
�@      @                �G���@      @     �5@�����?        �Y@�H��?                        XG��).�?                
3����      @                Q>��"�      @                w�{`j1 �      "@                ���mU���      @                w�{`j1 �      "@                ���mU���      @      9@r�H�d @        �k�g��?2��Y�S�?                �/�Ǝ?                ,�yo#�@      @                 "dO��@      @(�o|�Y�?�j�g���?        ��ݮ��?     �@@Z���r��?        ;ڼOqɠ?                ��X�櫿      4@                ��qT���      @                ����      &@                %������      "@                �.���@      @                I7%�/��?      @                �.���@      @                I7%�/��?      @                �#�����?       @                9� ��A@     �P@N���P�?Mp�@        b�/��?���Kq��? eN�Q@        ��Y@�H�?                "�v���      @                �����      @                O��@�     @W@                j�ȼ�a@      @                ��]��@      @                L��wO�      &@hyܝ��?c�럋,@              �?     �>@�6��N"@        ~�K�`�?      %@�Ӧ@        �h�>��?��N�`}�?nm?�^@        5�0��?      @��(�0X@        #Qj�a�?                a�;�<v��      :@                g^4��FB@     �R@                ����a�:�     �b@                �!q)�� �      ,@                ���vh��      @                ��!C0@      >@�.n���?��A�y�5@              �?     @G@"�{�@        ������?     �A@H��VJ@        mާ�d�?     �:@Dw3_�"@        �k�g��?      K@�(W\��?cA.eu?ֿ�k�g��?                �L�u�@C@     @T@                ���_�'�      9@                ��E`*�     �\@                (���@      @                |/v@\�*�      2@                ���<4�      K@��d���?�Q�nD:@              �?     �R@�*^���@        &C��6��?>�xM @���c	�@        mާ�d�?     �9@��Of���?        1��R�?                        ��ݮ��?     �V@*����+"@        �A�k��?Zd;�OE@�a�ANC@        {���?     `R@HE��oD@        w���L�?��#bJ��?�_N�K@        #Qj�a�?����?9�FQ$�@        Sc��|�?     �P@�1�J8�@        ��6�S\�?                j$����     @S@                X�׍"	�      "@                ��{��m-@      2@                �jQ���      @                ���;���?       @                ن�+�C�     �S@                ���;���?       @                ن�+�C�     �S@                �T�gD�      @                R3<�}	@      "@                .jc��G@     �T@                ��
)��      @.�o��%�?� ��:@              �?��s�/�?��ToqG	@        �۵r�3�?p=
ףh@���N�^@        �H�{��?                <�)�BC�     �g@                j�t5�      @`��"�L@`��@        �6�S\2�?Z�����?                �"Qj�a�?                HS�h-]�?      ,@                ǨL,uF@     �U@                ��Z9�;@     �L@                BH_i��0@     �E@���a��?�s�p��<@              �?ni5$�q�?�@��.@        �۵r��?��ʡ-@@S��O�@        @�H�{�?���v�? i��MU@        ��f�?      %@��9ȉ�@        mާ�d�?                �yg\�       @                ��q�xXH@     @Z@     �Q@��֬�@        i�>�%C�?                        )5�0ȗ?                �D�_���      @                {��-@      5@                �Ii��L�     �[@                б����      E@                �Ii��L�     �[@                б����      E@����y�?�V��T3@              �?z�ѩk�?<��}�@        �`mާ�?�z��{�?�����?        �>�%C��?�G�zO@%<�AJ@        J�=���?     �A@��Z���@        �g�t��?                �v��@      @                `<x��A@     �`@                ���G$�3�     �U@                [XG��@      4@                �T;cš:�     �G@                ��i�S@      @��a��@n���K&1@              �?Y���-�?����V�@        i�>�%C�?����1@���2��?        \2�h��?      @�¸���@        ��o���?�l�/�@�L����@        �H�{��?                ����'@     �E@                H�G��7@      E@                ��R�i�)�      V@                �^E�\�2�      ?@                $[C�R�(@     �T@                �m�)d�      *@�F ^ׯ�?(�oY8@              �?     @B@(��xC"@        �H�{��?���{��?�J���d@        �n��	��?      @BDD֔@        �۵r�3�?     �U@���7C�!@        ������?                ,� AN� @       @                P��=��=@     �W@                �g% ��@      @                Ǣ<�i��     �K@      -@]��y~@        }�(5�0�?     �Y@��H[S�?        �"Qj�a�?                ﾭlJ��      E@                �'��G�     �U@                N���j�?      @                qYQ���@      @^�,σ��?�_k��4@              �?     �:@|�)�W"@        ~�K�`�?f����@^K���@        �h�>��?      0@p��E3@        �D���?�ǘ��P�?���C��@        �0���?                ���ѱA@      W@                ���5���      @                1��Z�@      @                n����H�     �Z@                ���m�#�     �Q@                �y�$@      4@!Y�n�@0��p�6@              �?D�!T�Y�?켺�j9!@        �]+'<��?�T�t<f�?e��	���?        �D���Y�?                E����=J�      j@                ���Nn!@      4@                $��\*#@      @                n�c���:@      P@     �5@��,�@3@              �?      '@�R�k@        ��]+'�?     @M@�J���@        �"Qj��?     �G@�e��%�@        ާ�dֱ?|�͍��?�
w��@        �D���?                A���t2@     @X@                �N1(=@     �P@       @�%��@        p��Z9�?       @                ��ݮ��?Gɫs��?����@        ?�%C���?                        j�a�/�?      +@��ߤ8@        ��).��?��"��~�?                ;ڼOqɐ?                Г���*C�      Y@                �aFb�q@      @                9�����      <@                /[��\RB�      R@                ]4_&z@@�     @V@                �����S�      &@                        ;ڼOq�p?      B@i��.��@        )5�0ȧ?                �b�w ��?      @                T��C¸�      0@                �b�w ��?      @                T��C¸�      0@                s�p|� �      (@                p�LsK(�?      @��� ��?�����8@              �?�9#J{��?��oŏ@        �/���?      3@-Qᄣ@        �۵r��?�����?���_`�@        >��E��?cAJ��?L;O����?        )5�0ȧ?/�Xni�
@}�%@        p��Z9�?�5���@2|��zR�?        �Y@�H��?                5x֐CME�      f@                `o` �� �      (@                ��9\@      @                ��k��?      @                ���&��      2@                ��T+@      (@                �4P0��A@     @P@                ��h�L/��      @���[�?�. M5@              �?      X@b�_�d@        B�k�g�?�:�f�a
@��+q��?        }�(5�0�?      3@�c�T@        M�n���?��b('�?                ��ݮ��?                :���Q0@     �Q@                ���ܾk9@     �K@      @'a�;��@        �0���?j�t�F@,�	l�� @        f�"Q�?                2?er6�D�     �b@                LpT[f��?      0@                ��}��?      @                1ٕ�m�4�     �C@     �P@���hM@        UUUUUU�?l����J@붙Ԯs@        �v���L�?                W�D�9�      G@                �w�u���?      @     @A@qq$��@        ��ݮ��?^���T��?Ƥ�MM#@        ��).��?                ����&@      0@                ��5�dA��      &@.s�,&��?�s2È�@        �:ڼO�?fffff�N@E�1���?        ;ڼOqɠ?                䐅��      7@                �+d���#�      ,@                R �����?      @                %�S�b@      @��^�?�/&] <@              �?c�tv2x�?��X�#@        �0���?      #@��)R5@        ��o���?     �?@�g"HG@        �r�3��?                        �/�Ǝ?                �H����      @                PP�N�I@     �]@V�zNz_�? ��E
�@        ��ݮ�?      '@�0�p�@        ��:��?                �X�C$�F�     @Y@                �]欇��     �P@                �E�K�G�      X@                dΎl" @      @                ���ܹe�      O@                �[G��@      @B	3m�
�?�����k3@              �?     �6@�����g!@        ~�K�`�?b֋��(�?I+��*�@        �h�>��?0/�>:��?�QA�!q�?        �6�S\2�?pw�n�P�?n\qh<'@        mާ�d�?�MbXUh@,�\,@        �6�S\2�?                        XG��).�?                ̦�r�4�     �O@                m�B��4�     �@@     �=@�m̯��?        �:ڼO�?�0�*�?H$���@        �u�y��?                ��+p���?      B@                ��Sd-�     �J@���G��?���u�>�?        ��7�v��?                        j�a�/�?j�t��K@ ?py��?*[��)&�?��Rc�?                        j�a�/�?                �K���C@     �U@                �+�5/Z�      @                �Ͷ��@      *@                ��n�nB@     �R@                �Ͷ��@      *@                ��n�nB@     �R@                a�H�� @      @                �&�{��@      @                a�H�� @      @                �&�{��@      @f�c]�F�?)W+�C3@              �?      �?�,�I@        �}�K�`�?     �9@�g8?@        2�h�>�?2�}ƅ��?                ������?     �V@��D��o@        amާ��?                #PsCC@     �V@                ţ�;���      $@                �Zea�3<@     @Q@                ��w��@      @@                �ٗhv�H�     �e@                s�XG[�@      3@ o�ŏ�?k�Y�8@              �?      -@q��@        �6�S\2�?
ףp=zF@�w��x@        �!XG��?�q�Z|��?�\6@        ��!XG�?,g~5��?  GV�@        ;ڼOq��?                VM���      5@                R��C@     �W@                ��mh��      4@                ��W��@      &@h��b��?]��R@�U1пi�>�%C�?h��b��?                ;ڼOqɐ?                l�s�j�F�     ``@                d�*�      .@                l�s�j�F�     ``@                d�*�      .@������?Ч�&#s3@              �?�1�%$�?h���En@        Pq����?�=�
��?����?        amާ��?     �A@�&/@        ��|�(�?                        �/�Ǝ?                � T�/@      *@                ��޵
:@     �S@     �H@\"}�@        B�k�g�?     �G@����$|@        mާ�d�?                  pp�H�     `f@                /�"�ڜ@      7@                �q"f2K�     �d@                M��uX�@      ,@                ׽��S @      2@                ��c;3w��      @jo��ɔ@��5l�a*@              �?B��=�*@bV�	@        z��!X�?���� @�.EK��@        �:ڼO�?�x=�?�m��@        9����?                        �/�Ǝ?                Ζ���@@     �Q@                ��� ���      @                �3��@74�     �`@                �E2�,@     @U@                �3��@74�     �`@                �E2�,@     @U@O���|��?�m:��3@              �?D� ���?q����m@        [9���?��kC���?�����@        J�=���?���V��?�I.�*�@        ������?.�o����?                �k�g��?                �����D%@      .@                ;1�<�7@      X@                4(��X	C�     @e@                z$u� �      (@                ��z�bE�      f@                �|@-���      @��~�T��?�d6�+8@              �?^.�;1k�?34!�[
@        �S\2��?��1 {=�?UTHO�@        "XG��)�?                �*&l�'�      U@                ��9Y`�:�      N@     @A@`��`�'@        @�H�{�?���#b
�?w�)D�?        Z@�H��?                �|���      "@                ]�K�վ@       @                ���m�@      @                g���G@     �`@H��Q,7�?|�E��-4@              �?     @E@el�`�@        ���}�K�?     �Q@O �c6@        T\2�h�?     �V@�e�M!@        Nx��A��?     �L@�%��?        ^+'<���?                B�3�B@     @R@                j$�4�      *@                ��^XU_0�     �]@                ��� 7&@      3@                ��P�U�4�      C@                F
��!�     �B@��x�@��?n0�}�83@              �?hyܝu�?"�9ݍ@        ��7�v��?     �8@�x��L@        b�/��?                V����K>�     �Z@                ����XT�     �T@                "-}s�#@     �M@                �-_��;@      J@n��S�?�>+��#/@              �?      @�fx�m�"@        C��6�S�?;�f���?u��*��	@        z��!X�?     �3@w(g�έ@        j�a�/�?     �8@P����D@        }�(5�0�?                *W<�@      ?@                �CPt�BB@      S@                ��dq���      @                �:JD��"@       @      +@��[;@�d���8Ϳ0��f�?      8@��J���@        ��7�v��?                ��ܿ�8�      O@                �Ꭿ�+�     �W@      5@�u��T@        XG��).�?     �;@�l�X��?        #Qj�a�?                ��$�$��?      @                \$��      @                �P��N @       @                ����?      @n��S�?��;�6@              �?     �L@�6�8"�@        C��6�S�?Zd;�OE@'�K��\
@        z��!X�?                �@8JaD�     �e@                �����?@      @                m\�#���      *@                (�bA�OF@      [@���=�$�?7�of�1@              �?cE�ax�?dT�J��@        ��|�(5�?F�2Ɉ@���>��?        ��ݮ��?��&��O�?�d^#@        Pq����?                        j�a�/�?                �+O�ח"@      .@                ݲ����9@      U@                ��'Zg[B�     `g@                ����@      "@                ��'Zg[B�     `g@                ����@      "@MJA����?V�J�f/@              �?     �L@�3����@        ��:ڼ�?z�Cn�[@�������?        �y��!�?      @��i��@        \2�h��?^����?                XG��).�?                ����{%@      R@                �����?@      U@                "3��� @      @                �(���A�     �`@                �f&}�;�     �_@                H4��,�      &@���N��?�sl�1@              �?�����l3@�u��"@        - _$J��?j�t��K@Os�RsN@        ��A�k��?                        ��ݮ��?��Q��R@׸^ K@        8�v����?]����?�)k밖@        �}�K�`�?V-�M@�^�T\�?        �o��Z9�?                �� j�"�      .@                
���wC@     �U@                7�bD��E�      f@                �;@      1@                g+R6:�@      @                ��)P���      "@                �L���@      @                o�5PX6A@      T@���+�?�LU)A�-@              �?h��|?u�?�e	@        I�{��?`��"��>@ ou$;9@        o��	���?                �+>/�8�      W@                ��h��¿     �U@                [��3�
�      @                Zʲ��D@      ]@\�� �L�?��9B�~,@              �?��N�`}�?E u^��@        UUUUUU�?]P�2��@1�x��@        UUUUUU�?8��d���?+��}�!@        �k�g��?     �3@�ݦ�l�@        ��ݮ�?                ����G�*@      6@                &?��0@     @Q@      P@�m"� �@        �u�y���?,+MJA��?Td8�3�?        Sc��|�?                n
.�K�"�      "@                �u��ۿ      @     �I@�=w@        Qj�a��?     �P@ٚ���d@        ��E�Ը?                �c�sW�@      @                |����@      @                ���Z7�     ``@                w�v�?-�      9@     �7@                �"Qj�a�?     �R@�&�?��@        �]+'<�?                �@�Q-"@      8@                gD�w7��      @      "@�cG���?        �/�ƞ?      U@ ��F���?        �����?                �{|��ȿ      @                ��'4�      @                ʚ�x-t@      @                ��f'�	@      $@x]�`7��?�����/@              �?      @�X>��@        ��:ڼ�?�3K�4 @p=k4qz@        �y��!�?                        �/�Ǝ?      Y@*�d�(@        �/���?                Υ�8�U@      M@                �+/�t@@     �V@                Υ�8�U@      M@                �+/�t@@     �V@                Tb����B�      b@                2��2��@      @��m���?��`�L�)@              �?     �3@�6�t�%@        �a�/�?,e�X�@ ��@        '<�ߠ��?     �I@���ʄ"@        ;ڼOq��?     �=@�Ď�!�@        ^+'<���?                ���<j<@     �X@                R04֩
�      @      /@D/���@        &C��6�?      0@5��S��@        ��!XG�?                K
�H�     �X@                q�ݟ�C�     �K@                �v@      &@                l�ʊ5�      ,@                �A���      @                wk[��+@      &@�q�@H��?�""!^6@              �?fffffT@̬+�!@        ;ڼOq��?u�����?!(�E@        �K�`m�?+j0��?&�����@        ��	��7�?                        j�a�/�?                (�2�Ү@      @                �}$�6D@      a@                ��J@�     �a@                ����Q�!�      *@                ��J@�     �a@                ����Q�!�      *@>
ףpeD@�=�-�(@              �?��MbA@���^U1 @        #Qj�a�?"�*��|�?[/p@        o��	���?                N��&�     �H@                �{F���-�      :@                ��w�,!�      R@                n�9�'B@      c@֋��hw @����X,+@              �?h��|?u�?Z�9��@        '<�ߠ��?�r.�5@s��)3�?        ��Y@�H�?      @(����@        b�/��?      *@y�7s� @        �a�/�?                ����@      $@                ��!Ƥ�7@      V@ףp=
E@-��-@        XG��).�?����?ǽ�=%@        �a�/�?#�-�R\�?Y�Z�l�@        �/���?�mnLO�?�`D���@        �g�t��?                �8���
�     �H@                &�}�Y�'�      4@                ZG�җ<(@      *@                O$j����      *@                �2EF�n@      @                x?R1���?      @                ���ܢ@�      T@                r�<E��?      1@��~j�$G@J��h�o&@              �?�����l3@j _��/@        �����?p���T��?�J��q�@        �).�u�?                BA_#��@       @                �#og<�     �W@     �C@����f�&@        s�3���?0�AC���?��VMk	@        �r�3��?     @@@M�t
�0@        ��o��?      >@��=�.�@        i�>�%C�?                I�~LWA/@      8@                �a'�.:@     @Z@                �N�U�N,@      6@                :ۣ�2�
�      @                ��`�>p3�      ?@                v�Uq�?      "@׆�q�&�?�R��!@              �?     �2@�{X|-@        C��6�S�?���ׁs�?/V���?        z��!X�?     �X@�*�$@        ��Rc�?      #@O<��ӳ@E{�����0���?                /FT��@      @                ���k�3@     �Z@                �,���1�     �`@                6/=��&@      0@                ��FS�@      @                t�$���5�      A@1�Z�H@]f��6-@              �?     �:@[?U �$@        7�S\2�?{�G�>R@�CK�|@        e���}�?Ǻ����?���w@        ��o��Z�?     @A@�Ի�@        �Y@�H��?                `���0@     �^@                ؄�Ӵe3@     �H@l�����?)�S���@        ��L�n�?�(\��%C@J���ڷ�?        �/�ƞ?                T�� @      @                �g� ��?      @     �R@�x�*�@        �h�>��?�ʡE��@@!�4��?        �Y@�H��?                $z�N��?      @                �w@+@�@      @ Ϡ��@�Ip�(w@        ��Y@�H�?      0@RwAR@        )5�0ȗ?                 Ⰺ��      @                ORg��M�      @      C@�f,�v�?        �Oq���?                        ��ݮ��?                        XG��).�?                        �"Qj�a�?                z���wQ7�      D@                �����1�     �J@                z���wQ7�      D@                �����1�     �J@                z���wQ7�      D@                �����1�     �J@                z���wQ7�      D@                �����1�     �J@��ek��?P��R�%@              �?     �6@�x����#@        ܵr�3��?)\���Pc@��q)��@        I�{��?      @����@        p��Z9��?     �F@�&��M@        �n��	�?     �K@����\�@        ��}�K��?�(\���@|�5��"@        �k�g��?                        ��ݮ��?      D@�O}�r��?        ��L�n�?     �9@�
"�k(@        �y��!�?>����,�?r�F�y
@        +'<�ߠ�?                �t����=@     �R@                T���kd��      @                        ;ڼOqɐ?�G�z�e@���P#��?        ��ݮ��?                ���g�      @                Z��?@      &@                I[QP��      @                ��g���	@       @     �0@+���� @        >��E��?      G@=KZ<��@        +'<�ߠ�?                2��:|�,�      <@                ����#�?      @      ?@�ɗ��[�?        ;ڼOqɐ?     �C@�w�@r���?�0���?      H@��{@        ��|�(5�?o*Ral!�?�L~L@        ��ݮ�?                ��h+z��      @                ����eA߿      @     �;@��\R�&@        #Qj�a�?     �7@,2��I?@        ������?�Y��B3�?                �"Qj�a�?     �<@��՚�@        ������?                �0/��3@      1@                J�q�t@      "@                �0/��3@      1@                J�q�t@      "@                ��8G+>�     �F@                �W�Ò~�      @                �x01��:�     �G@                �6	���      @                �j��@      @                �a�qj�?      "@     �8@�
�9��@        ��Y@�H�?                        �/�Ǝ?�䠄Y�?                ��ݮ��?     �K@�?����@        )5�0ȗ?L7�A`e�?�2�,�@        j�a�/�?                        ;ڼOqɐ?                x���uk6�      D@                �M�֪@      @                i z��4�      D@                �HrE5��?      @                        XG��).�?                        �"Qj�a�?���kq�?��Lœ\�?        ;ڼOq��?                        �"Qj�a�?                ���Wj^8�      B@                ,Wt�J/�?      @                ��[��4�      @@                Z���"�      @                ��[��4�      @@                Z���"�      @                ��[��4�      @@                Z���"�      @                ��[��4�      @@                Z���"�      @)?�����?�����!3@              �?     `b@9$�\�'@        E���Y@�?��1ZG�?$\���?        w���L�?V-��F@�F��'@        '<�ߠ��?��Q����?                XG��).�?                �J�AT	@      @                Z��1�<@     @U@                �Wb�#hF�     �U@                �1gX�3
�     �]@                �q#��cD�     �h@                ��*�U;�       @_�L�j@*5�M(@              �?     `b@z�u�w&@        ��	��7�?�G�z^E@m��	�@        ����, �?      @fDr"@        Qj�a��?s�FZ*��?4-�fF��?        ������?                !V�����      @                ��%Ç<@     @R@                        ;ڼOqɀ?     �<@[�:c.?@4ʞsх��v���L�?                4�ǯ@      @                ���c�@      @                4�ǯ@      @                ���c�@      @                b�
�1A�     �X@                	ø����      [@GɫsL�?]ԕ6ZK%@              �?8�9@p�?��o�Z�@        �E�����?���S�%�?��O�f@        t�VNx�?                A�� Rp�     �f@                [oTx��       @                |xB@�<�      @                ͎�l�C@     @Z@��jHܣ�?mG25n�.@              �?��I�r�?/K(��@        �h�>��?     �=@�Te%�@        �).�u�?                ��!~�C�     �f@                #מ�v@      $@                }���1A@     �Y@                B�ю��      @0L�
Fe�?X�T|+@              �?     �:@G��δ�@        mާ�d�?���Y@k�:�d>@        ������?     �<@�Ԙ@        ��|�(5�?      >@a��KV@        '<�ߠ��?                0&m�S+@      ^@                �)�S5=@     �T@                [�LJ!�     �@@                �O�q�!@      .@                ��UF�Y8�     �E@                ���f#��?      @�1��o�?w&���4@              �?0��{���?���)@        ��f�?��jeb@��컆@        ܵr�3��?82���@�?�3���@        ��:ڼ�?]��k�?I�Qz�?        j�a�/�?                w�p��,@      W@                Y˻�G*6@      J@                P��:��>�      U@                �̷O��      N@                ��l���      @                �&;�g�      @���x�?է�|��*@              �?0�[w�T�?��"�P@        Pq����?�'�$�@"@����?        amާ��?     �X@#x��@        {���?�Fw;S�?�[Vm��?        Sc��|�?                 ƄG��&@      5@                ��h=Xk,@     @P@                =<e��H�      g@                ��:��"@      3@                ���?�k@      @                ب�E�@      @0i��Q��?������%@              �?ƊL���?�* ���@        amާ��?^��K�??�0�@        ?�%C���?                �[5���@�     �e@                ��@X@      *@                �˫z@@     �Z@                �a�ײ��      @uv28J�?�4���'@              �?     �=@j�=o��@        B�k�g�?� �> ��?�gǴ@        _$J�=��?     �7@�V��8@        �ߠ۵r�?BB��?�=�s�@        �]+'<ӿ?                ����M@      "@                W	x���>@     �d@                �֩��<&�     �J@                *K�Ģ�@      B@                >�/�)2�      >@                ��v��9�?      @��	my�?�����&@              �?      @5�]���,@        ���}�K�?ĔH���@�-;��?        T\2�h�?      3@	��q�?        ��ݮ��?     �Y@���$@        �a�/�?                z�����#@      3@                `L�6s1@     �Q@                �k��@      @                �i03Zb@      @                ����F�      f@                �>ˏ%@      7@r�t����?�+KE��!@              �?N^��?�d��A@        E���Y@�?:ѮBʏ�?\���Tf@        ^+'<���?                Z*�k�:�     `b@                �	�_�@      "@                _�,�U~@      $@                ��H��7@     �`@
ףp=zF@c��/&@              �?      '@i���$�#@        �/���?�� �rX@@,���?�#@        8�v����?      @��y��@        w���L�?      /@�į�`�?        ������?                ��I4�"@      @                #?��j4@     �f@                ���#�@      @                ��Κ%!C�     @W@                vB	��@      "@                o�$�?      @      #@����o#@              �?     @Z@}DvFH�@        ~�K�`�?��H.���?EwTM;�@        �:ڼOq�?      C@��/@        e���}�?      -@DV���@        ������?                �Qz��      K@                �Bԕ��C@     @^@                !�U<h�     �M@                �~��:6�     �L@                ��!Z��?      @                ���2�@      @�I�5�/�?��/6(@              �?     �C@g2~X@        >��E��?��Z��W�?yG��s@        �g�t��?                \�GFB�     @g@                k.��-@      1@                �2 �^�      "@                g��Q��?@     �U@���a��?(B}��~!@              �?v�ꭁm�?�A@�1@        �۵r��?       @Ǜ��7�@        @�H�{�?Է�鲘�?��5,F@        �r�3��?��\����?�ۺ^Q�?        ��!XG�?                        �"Qj�a�?      %@6돕��?        )5�0��?                ��n�,B�      @                ቮ���8@      \@                �4MY�@      0@                �JaD1�0@      X@��y���?��粵@        �D����?                        ;ڼOqɐ?                �!~�R�      @                �hU�r�      @                c�+�1'�     `b@                �LÁx,�      6@                c�+�1'�     `b@                �LÁx,�      6@���~�z�?Vg��:�-@              �?�M(D�a�?�[��lE@        ��:��? R�8���?�>�P�?        ���}�K�?��Hh���?Ye�PF8@        ��]+'�?     �@@'�n1�I�?        �"Qj�a�?                ��h�,@      9@                1	c��3@     �S@                ���K=�     `f@                2�Ł�@      "@                P��%��      @                _�#.%�      @���?�r^�ˬ&@              �?      @J�Py�� @        1��R�?      @|rL�U@        ��o��Z�?     �>@Ě@�K��?        ;ڼOqɠ?      +@
u�B@        �=��E�?                ��E�JU@      "@                S�J:M4@     @[@                �;1�q�?      @                �	���@      @���B��?Z!��%�@        ���:�?     �8@11���]@        ��L�n�?                ��_��>�      L@                i_n��?      @                *��A�(�      X@                Δ���@      0@      #@!n�Lk&@              �?�l����H@���t�@        ~�K�`�?      )@X@���@        �:ڼOq�?                �Rq��>�     @T@                ���J@     �G@                �`��@     �R@                ��.��;@     @X@˄_��M�?( I�#)@              �?      -@��E@!�@        h�t�V�?��N]��@��9�~�@        1��R�?                ?����� @      =@                R��c�@E�     `f@                }nŮ@t*@      8@                �Y��@�(@     �P@      @M�}d@              �?      �?���^�a�?        ��Y@�H�?     �5@w[$�"�@        �g�t��?                p/�h�u@      @                ���_@      @     �8@6���:!@        ���Y@��?     �D@���d&!@        �k�g��?
3m�ʊ�?<����@�m��;�пL�`m��?     �<@��ٞ@        �]+'<�?�P��C��?^�
��B@        ��|�(�?�e�I)(�?G]˞�@        ��!XG�?                z��8:H3�      Z@                �%��+;,�      0@                b�b�I	�      &@                }v��,@     �D@                0 /O� �      N@                M����q-@     �C@                �W]��'@      "@                �H�#�@      "@�wE�U�?�70��'@              �?      X@���5�!@        >��E��?�7�06�?�aYy:�@        �g�t��?                #^k�<�     `g@                K����p @      $@                +W���LA@     �X@                ���� �      @5^�I:G@SFb�'@              �?     �X@-U��5 @        4��]+�?ʉvR~�?���  @        f�"Qj�?                S��1<�     �Y@                ����/�@      @      @JҾ�7�@        �n��	��?D�l��iN@3y��;
@        �K�`m�?                Nj� ��@      @                ���|p'�      D@                s�A�q�:@     �J@                ��է}2@     �W@!Y�n�@�d+q�R%@              �?     �8@��<a�3@        �]+'<��?�����@�bu�K��?        �D���Y�?                ���^.$@�     @^@                �d���0!@     @X@                �5
��*@      >@                E5֔�J(@     �I@N�St$�?������0@              �?      @����T$@        ��Rc�?��C�lG@;��@        �t�VN�?      @A�O�j� @        �k�g��?�����<@�ÿ��@        Pq����?@�z��;�?J��I\@        [9���?0�AC���?)��n$�@��»�?��o��Z�?                \E҈�@      @                �k㤀�?      @                2H>O��@      $@                +w
0�]G�     �^@                K��� �"�      1@                B�_k�d@      *@                �n��,@      6@                ���;O1;@      Z@�vö��?%��)��#@              �?     �@@�WݤD,%@        ��7�v��?{�ᯉ�?��;�0�?        b�/��?      @iL�ª�@        ݮ���?     �>@U�Ax
@        @�H�{�?                =>O�h�@      @                O�Σ_7@      X@                �[��f@      @                D]oY^B�     @d@                �aS���*@      .@                $����-ۿ      ,@��{��D�?�*� �m'@              �?(I�L���?w�#M��@        $J�=��?[rP���?� ���@        �k�g��?                 p�E5�     �d@                �R�@Ҷ�      @                        XG��).�?)yu���?e!���@        }�(5�0�?                ��6w�
@      @                ���N%�:@     �^@tA}˜��?F��S��@        ާ�dֱ?~W�[��?oZ q� @        �g�t��?      C@�VU\�@        p��Z9�?                        ��ݮ��?                �ݝ��V'@      5@                �@�1@     �U@                �HW���@      @                ���J�      @                �HW���@      @                ���J�      @d�����?->���.@              �?     �1@]�_|��!@        ��o��Z�?�����?qĕ�a @        �, _$J�?*���P�?#�Dt7��?        ��6�S\�?     �6@#��|�	@        �D���Y�?                ,i�8J^	@      @                ��@@      b@                W���<�     �Q@                �;�<kC�      "@     �2@��Sʕ�@        ���:�?     �8@�N���]
@        ��ݮ��?                �{�v���      "@                ��du�$@      5@      -@�3V)(��?        ��Y@�H�?���N��?A7�+۹"@        [9���?                �6��      @                �tV�G�      @                ZO�Z��      6@                �=�B)�@      "@���EA @��<��� @              �?      @�1Θ1m@        ��ݮ�?B��=�*@C*'d7�?        >��E��?                        �"Qj�a�?     �>@��-[@        UUUUUU�?                �[�dL@      $@                �ʈ��$1@     @X@                �[�dL@      $@                �ʈ��$1@     @X@0�*���?S��@        �	��7��?     @H@�w�qT@        �۵r��?                ���u�9�     �Y@                z;�$ �      $@                �{5e "@     �K@                ���^�      5@��k�U�?��j�.@              �?     �3@�k�F�@        Nx��A��?�<I�f��?����ȏ
@        ��, _$�?      '@,������?        2�h�>�?     �6@���1 @        p��Z9�?     �6@                XG��).�?�)t^c7 @�S��\@        ��o��Z�?                jƍ� !�      8@                �{��A�      U@                ���%@      4@                �&����      $@                ���%@      4@                �&����      $@                HY�xa�޿     �O@                �%�}6@      W@(\���Q@���b��!@              �?     �V@��� �p&@        ��:ڼ�?8�A`�@X@_����?        ��}�K��?
ףp=zF@TI��gu@        ���, _�?�G�z4A@[ê��@        ��o��?                ��;�5@     �G@                "�5�j�@      7@���Q�C@�j���?        &C��6��?     �R@v���@        �n��	��?      .@ =��m�?        ;ڼOqɐ?     �8@1H�2"@        �g�t��?                ��aR9�-�      S@                �?z	�f(�      8@#��~j�K@c�i��5@        <�ߠ۵�?�����J@D_�J��?        ;ڼOqɠ?                ^F�-�&@      F@                s\��@��      E@                ��|�2�      @                )B�a�"�      @                T�4t��@      @                J;����@      @     @[@|1��1�?        ��ݮ��?      1@�Q�˺�@        p��Z9�?                �`����      @                ����>p�      @                eG�mq��      @                i�]b�'@      (@b�� � @4�.q�L!@              �?     �8@�([�{@        
��7�v�?^��K�?ؤ�)�@        �a�/�?     �2@�c4��@        G��).�?     �\@A���@        ��E���?���Q@@)�'�@        �Oq���?���	.� @r4��V�@        �"Qj�a�?                dU��Z��     �B@                �#�P%-@      F@                *�gOU�>�     @[@                �����@      "@                ��6�"��      @                �%���@@     �V@                        �"Qj�av?                        ;ڼOqɐ?                ��>}���      @                Hk処0�?      @                ��>}���      @                Hk処0�?      @��Q�-R@hA�iD�"@              �?ʡE���E@�@�@        Sc��|�?ףp=
WA@s��#p�@        �r�3��?                ��q�(�9�     �Y@                �q}�@     @a@                �>5�2@      @                㫾ɐ�/@     �K@r��]��?=�jG�M(@              �?z�ѩk�?�+i�@        �����? �	���?�~�_��?        �d����?     �;@��ȁѰ@        J�=���?��<�;��?Cő�� @        �t�VN�?                .�����@      @                ��3�3@@     �`@                �y˩v$@     �P@                ~ �z])�      A@                �4��jm8�      L@                ����8q@      @fffff��?K�6�M� @              �?0��{���?䢯��u	@        ��o��Z�? <�n�?aT��@        �, _$J�?S��.��?p��	�@        ��:ڼ�?Բ��Hh�?��
#s@        )5�0ȧ?,�)��?ø����?        )5�0ȗ?*:���?�tQyUa@        q�����?                ��/i�@      @                �憃#�@      @Жs)���?F��Kb@        �/�Ʈ?     �2@���v*@        o��	���?��� �6�?b_8�a@        #Qj�a�?J�i�W�?��
X�?        �}�K�`�?                ['g'!S�      @                ����!>@      ^@                        XG��).�?                        ��ݮ��?                 	����      @                �>Uӣ��      @                 	����      @                �>Uӣ��      @                 	����      @                �>Uӣ��      @t^c����?VY5�)@        ���}��?|�/L�
�?�5�@        ;ڼOqɰ?                �����?"�      (@                `ɐG~��?      @                Yh�:U��     @V@                �Q;�7'�      ;@                �!�@       @                ��G\��?      @��ek}��?�tVi� @              �?     �F@z1�f� @        8�v����?|�w�@{��3	@        �/���?     �8@�1մ��"@        �(5�0�?     �H@��n�@        ާ�d��?                !�9�=@      [@                ���N-S�      @      @�R;��@        �"Qj�a�?�����?                �Y@�H��?                �`���,)@      <@                =|;���     �M@                �@VT�
@      @                YV����C�     �V@                �Hv�9*<�     �S@                ���z�<�      .@��~�T��?��>�@              �?A�c�]��?vD
�u@        ��, _$�?      /@@����Q	@        ��L�n�?                ��fB��     �l@                �E�].C�      &@     �5@L8��P��?        UUUUUU�?                        ;ڼOqɐ?                .�8���@      @                �F��2@      J@                .�8���@      @                �F��2@      J@      @�A(��L @              �?      �?��`�{Q�?        +'<�ߠ�?b�� ���?K��n�#@        {���?                rj8p��@      @                 d]_'%@      7@      @����3@        Z@�H��?��(\�jh@�����k@        �u�y���?�)�D/��?�����@        ��ݮ��?      !@Zc-Jg��?�_-Ҙ��e���}�?�]P�2�?��L,N�?        ާ�d��?�o|�%�?�$v���@        ;ڼOqɐ?                � �S��@      @                �F�V��?      @                � �
>�5�     �P@                j2R��*�     @\@                ��'�ĳ
@      @                B�?N5@     �R@                        ;ڼOq�p?                        XG��).�?                rw��4��      @                �����?      @                rw��4��      @                �����?      @     @Z@�G4Jk'@              �?��x�@������+@        [9���?l[�� ��?�u�n@        )5�0ȷ?���)Q@`ɣ� @θc����H�{��?�G�z^E@TC��� @        s�3���?                        �k�g��?��n�?�/t�~[@        ;ڼOqɰ?     @G@tդ9@        ��:��?                        )5�0ȗ?                ����]�      "@                �/��@�6@     �Q@                ����]�      "@                �/��@�6@     �Q@     �_@��?        �}�K�`�?j�t��@t
x&h�?        �u�y��?      @.��]�p@        0��f�?       @��2�@        +'<�ߠ�?                ��#��BG�     `d@                �{�XO@      ;@N֨�h4�? ��K@        #Qj�a�? <�n�?\��-�?�:pY�ÿmާ�d�?                        �"Qj�a�?      R@������?        ��E�Ը?                        �k�g��?N-[���?                j�a�/�?                1{#�VA�     @_@                5��z��.�      <@                1{#�VA�     @_@                5��z��.�      <@                ��MI�gE�      b@                �2U�1�      "@                ��MI�gE�      b@                �2U�1�      "@                d+�j?}@      0@                IX6ƭw@       @                ���f�@      @                �i��q�@      @                �"7�</@      @                *�y{u�?      @z�G��?���\M!@              �?     �8@��uà@        �d����?�ME*�-�?��[\%$@        �6�S\2�?     �@@�����@        ڼOq��?82���@�?�F�]�@        �}�K�`�?                $�PƲ@      @                ~��,�08@     @W@                ��r�p�@�      d@                �����X"@      9@                �E���O��      @                ���P-6'@      (@     �2@P�<��"@              �?      )@k��j�@        ��7�v��?     �A@���XR@        ��D��?                        XG��).�?     �A@5��@        �{���?J+�&@@<��v@�G�?�?��ݮ��?     �Q@(Q�m�@        �D����?                ք^CA?5@      J@                8U����?     �[@                ��ЈG�     @P@                ��'�T	=�      Q@                ^8ޞ��      @                ��%��7@     �F@                ���sw�      S@                 =H<P @     �A@��Q�I@[�5s�&@              �?      -@~ ��3�@        �{���?     @O@�"Vj@        �r�3��?                YtՋɩB�     �Y@                IZiDa@      ;@                �k���?@     �\@                )�^%Zv�      K@]��+�?\���D_!@              �?ҩ+����?p�N�@        ��o���?���P1N�?�>X��Q@        �0���?     �B@,UEp�$@        �6�S\2�?      #@0�2�@        ��o��?                Ȣ�bu�@      @                �ȇ�k4@     @d@      @�j���X@        ާ�d��?      F@$��K�@        �u�y��?                �����u1�      =@                �U��^X�?      @                RD�z�
@      @                	�K�5�      U@                w�,���?      @                /�*�W @      @�P�fo @���x|@              �?     @O@1}*�R@        4��]+�?�&p�@�h�/e�?        ��D��?                �5��3+8�     �d@                �OH)@      G@                >0���.@      A@                {oug�`"@     �K@L�ԲU @! ��l @              �?l	��gs�?�ī9Gp@        �h�>��?�!�uq;@@�����?        �).�u�?                ��4�'�     �d@                p��s��.�      C@                �+<@     �I@                @�E��.@      F@0�*��?}�;�c�%@              �?     �R@���F�^%@        ��Y@�H�?2���s�?_2M��?        ��L�n�?Жs)���?^��N:h@        �0���?     �T@`�8{~��?        �k�g��?                !-y�M@      @                *�OY k5@     �X@                �����%�     @[@                H�|_7=�     �P@                ƶ��p�@      @                ���:@      ,@��x�@��?�G��+'@              �?�;����?������@        ��7�v��?     �=@܌f�e@        b�/��?��@��G�?�<�=�@        �۵r��?                        �}�K�`�?�٬�\ @�j�����?        ��ݮ�?                        �/�Ǝ?                bV4�"@      2@                .�}�m3@     @S@                bV4�"@      2@                .�}�m3@     @S@      �?��u6��@        $J�=��?����9��?"��ɦ�@        �k�g��?                ��\��e?�     �f@                �ʠqv@      ,@                        ������?[rP�?ĳ8�K+�?        ��o��Z�?�ek}���?K{)����?        �u�y��?                        j�a�/�?                "o�@      "@                �]���k��      @                $LL��1?�      e@                ����x��      @                0|��q@      @                �$�Yx�@      @                0|��q@      @                �$�Yx�@      @HG����?+��"R"@              �?     �:@��G�@        "XG��)�?��#0�?��+SSq@        �Oq���?      @������@        amާ��?      '@�#Kp�@        �����?                wB���@      @                ����0@     �U@                ��,�!
@      @                ����D�     �g@                `�m�O�@      @                ���yx���      @fffff�G@*h4���#@              �?      H@R�R@q"@        �`mާ�?l����J@�7��;�@        �Oq���?�G�zN<@���9�@        WNx��A�?���Q@@�_ɗ���?        �"Qj�a�?                �·�3�3@     �F@                ��4u�;@     �b@      @c��@        UUUUUU�?J+�&@@(��eW@        �"Qj��?                QZ���Y�?      @                �-��eQ@      @                a�B���?      @                H��k-�      9@                	��@       @                ��}�s�&�      O@���=�$�?>
��O#@              �?"���?�@���#@        ��|�(5�?\*��{@g�e�p�@        ��ݮ��?��jH�c�?ڂ��8@�E�6N䴿�۵r�3�?�x]�?���af��?        #Qj�a�?                �49O�=@     �W@                ��疀��      @                ^�A]�9�     `g@                �ڇpY�      @                �O��@      @                ���� @      @��ek=�?Q����$@              �?�L��;�?BN�ty@        ��:��?ı.n�A�?Fv�]��?        ���}�K�?                ��s�~�6�      h@                V"yq�n�      @                ��8��@      @                Jt�M�4@     @W@[|
����?\���w@              �?�,	PS��?v�r��h@        _$J�=��?��:�q�?~��M5�@        B�k�g�?F��_��?�H�@        �d����?����7�?|�c@        �/�ƾ?                �ՅIf�)@      7@                ËȄ�^2@     @Y@     �D@9�Q@        �E�����?                        j�a�/�?                ��'Y)�      :@                ��]I�?@      @     �A@�<S���
@        �����?     �:@��[�� @        �g�t��?                 L��B1�     @Z@                �Sw�q�(@     �A@                �X@2q&!�     �V@                ]�W�&_!�      ,@                0��6:�      &@                ��v�z0@      8@���)���?-r�F�%@              �?�(\��@�=����@        �|�(5��?GɫsH�?މ��@        ��]+'�?��ڊ�e�?�D�-��@��@���Ŀ�K�`m�?���6���?�.;lo��?        ��Y@�H�?+~����?l��Aʶ?        ��ݮ��?J�8��% @8V�UX�?        *.�u��?���9$�?��r7@        ��6�S\�?� �	��?�3d�@        i�>�%C�?                ����!B@      &@                ����@      ,@                (�y��@      @                �T^Y�
@      @                FJ��..@     �L@                �H�U=��      @     @O@u�2j@        �(5�0�?      #@��~D�i"@        ��o��Z�?                ���iOʿ      $@                ��ɦ�<1�      <@                0�ҹ�<�     @Y@                I�AR�
@      @     �1@omM��@        �y��!�?      <@o"��ż@        �Y@�H��?                        �"Qj�a�?�	���[�?���m�?        UUUUUU�?     �6@a��71&�?        j�a�/�?      U@n(�d�G@        mާ�d�?                /�o���#@       @                ME��;�@      5@                ��+"���      @                n
83Ļ(�      7@                ���	Gs	@      @                o��q�e@      @                V"�ۑW�      1@                ���-�@      @     �8@ZA)�3@              �?�Hm��?�H_�s�@        �, _$J�?     �;@,��u@        x��A�k�?d�`TRg�?��u秂@        5�0��?���9�?��Q��?        ;ڼOq��?                �5�i3@      A@                �	E��@     �O@     �>@���	6@        �`mާ�?                        �k�g��?                �|x�@      @                D�S��@     �A@     �D@�Q�q��@        s�3���?     �S@�=���@        p��Z9��?                FH�m�O @      ?@                WX6��<�     �_@                �_ݑ�@      9@                 ����@      @                �%!��9?�     �\@                -jV��@      &@��mnL�?�\��E�@              �?��++M��?�x
^@        �u�y���?��&N�@�����?�?        �).�u�?     �Y@T�RO�@        ��6�S\�?                        ;ڼOqɐ?                ��횻'@      $@                LҪ=��"@     �@@                �5.�<�     �l@                T��ص�%@      8@                �5.�<�     �l@                T��ص�%@      8@X��jN�?yy��$@              �?     �@@[��M^@        >��E��?%��C�A@�X5/@        �g�t��?����?�9K�E@        v�y���?     �6@Ϛ� �<@        @�H�{�?hDio��?��(�ZV�?        ��ݮ��?<�O���i@����B@        ��).��?�kC�8�?������@��8L����(5�0�?��(\��A@��K�!@        @�H�{�?     �7@SX7�:@        @�H�{�?     �8@��1��?        @�H�{�?                �ߦ^�j�      @                5���;�
�      @                n�v��@@     �W@                ��M�.� �      @                �r�vʰ�?      @                ��."@      @                h�~B�      @                K���,�?      @                I���{B�     �b@                h����      @                        ;ڼOq�p?�Q�Q��?tx]A?U�?        �"Qj�a�?                ` �4f��      @                ��	xF� @      *@                r9��@      @                T��sq	@       @     �<@�:L_ʻ@              �?     @Z@����I�@        mާ�d�?      @�}ֱ��@        �K�`m�?                ��%-�     �k@                �	��ET�      @                �Z�_�+�      "@                
�N@f�6@      P@      (@>�)��t@              �?                        �k�g�{?     �2@h�%� @        )5�0��?                nH��l@      @                6�]��T*�     �r@      B@�/���}@        #Qj�a�?     �:@M*v͒�@        �/���?                ��A����      (@                V�Ң2�      @     �7@�].��E�?        &C��6�?      +@{�0�4@        ��Y@�H�?                ��PD�*@      &@                ��&�p@      $@      @�4��9&@X˶m߂��^+'<���?     @Z@��)Ie�@        ��d���?                StmG�@      B@                Q��|?c@�     �^@�/�$F�?�=ҭ��@        ������?     �^@��Ƌ7��?        �}�K�`�?     �P@�b��j @        ��).��?      0@@��%i��?lwmcܧ?�).�u�?                ��O@      @                "5�<@      @                z�#�w3��     �B@                �J����      "@                �L���U�?      "@                ]�,�5�+@     �B@�?ޫV��?mIBs@              �?�U��y$�?U|+���@        �VNx���?n��R�?.KZ�@        ��f�?      -@���1�@        ��E���?     �F@bK��D�?        �}�K�`�?                #����� �      @                ���z�2@      O@      )@�z���@        ާ�d��?      @"�`@        ���, _�?                Z@��	�      @                ��;	��      @                ������      8@                <����M-@      5@                c�H@      @                �-Ŋ!B�     `f@�E���$F@z�� @              �?      0@��z@        2�h�>�?     �O@�����@        �}�K�`�?                <���:�     @R@                �r�|�@      ;@                �M��q@@     �g@                �PQz��      $@9{ڡ�?>@oqW(@              �?     �Y@�f�u @        
��7�v�?���B���?���@        �a�/�?x�W�L@j�U��;@        ��ݮ��?      _@������	@        �ݮ��?                O�u%:@      @                {�����6@      W@                c��{IC�     `e@                ������@      (@                ����_.!@      "@                ,`&���?       @dX��G�?y�2
�@              �?     �:@�2�g�>@        �0���?�CQ�O$�?��c��?        ��o���?      -@jܠ�Z@        �D����?      C@��^���	@        #Qj�a�?                ��(%�@      @                �r~�-@      ]@                h��v:�     �U@                w;�����     �T@                 �Ƹf��?      @                v�F�@      @���?�M%�A@              �?      @��/��k@        1��R�?:��H��?���t�[@        ��o��Z�?                @Y`@       @                �����;�      f@                ��@�1@      A@                ,��x�@     @T@      '@#�ط�@              �?      %@v�'��Y@        ��ݮ��?Z�!�[=�?�3�2̘@        Z@�H��?                ;bK5�@      @                �����s!@      C@     �S@@</ @        ��|�(�?�P�f�@.�w��@        )5�0��?                �Zu��I?�      h@                �Vҡp;@      (@                �Mp_#-@     �C@                `����N �      *@�Pk���?zB���]!@              �?      -@&^��
@        l�g��?      ,@ͮ_m��@        J�=���?                b��7�1�     �D@                G�Tt��      L@                A���     @^@                I0�`��>@     @T@ �4��?d��d�M(@              �?��9̗W�?�Q2��i
@        ��|�(�?��+e�@)E���@        ��ݮ�?     �A@ר���@        amާ��?                        �k�g��?                B�˂@:@      Y@                l�3a0�      @                ��}�D�     `e@                gm�C @      2@                ��}�D�     `e@                gm�C @      2@��~�T��?�D|G@              �?H�z�;@	�#�*W@        ��, _$�?     �`@�px0�	@        ��L�n�?ffffff4@�Bb j�@        �f�"�?�� �r�a@d�̳6,@              �?                �?��Z51@     �K@                e�x����      @                ���ʿ      "@                k�v6A}#@      (@                {=���5@�     �j@                >���      @��&SE�?ha��qX @              �?     �U@RrZ��x@        �}�K�`�?��� �?Ҋ�Q}�@        2�h�>�?     �O@�����@        ������?     �0@>3��Y�?        XG��).�?                �G� x+@      ;@                )�.Ȋ�,@     �W@     @@@�;���@        �ߠ۵r�?     �4@��&��?        �f�"�?                7I-�,p�?      @                �>�R@      @                6���)� �     �`@                ��s�T&�      3@                �n9��K�?      @                �@�ǯ&�      0@@���,�?S�v�`&@              �?     �E@�{���'@        ���Y@��?Qk�w���?�K|�n@        [9���?      @����@        t�VNx��?ZGUD�?����7�?        Sc��|�?                        ��ݮ��?6�;N��@���i��?        q�����?                        ;ڼOqɐ?�ڊ�e��?�\����?        ����, �?                �(>��@      $@                {�獠�?      @                �(>��@      $@                {�獠�?      @                ���O��@�     �i@                 �����      @                ���O��@�     �i@                 �����      @                J�ʆ|
@      2@                ,�iB��(@     �G@     �]@���Q3@              �?      ,@dRR��@        mާ�d�?     `b@G$�\��?        .�u�y�?                W�",A�     @e@                �jL�,�)@     �Z@                l�X��@      (@                <tC;�@      $@     �X@���_��@              �?      /@r~�M�> @        f�"Qj�?     �\@7�`�}�?        ��7�v��?�,C���?�U��@        j�a�/�?     �<@�.��ͷ@        ��!XG�?                �����@      &@                LD[%W@      ;@                \�9
{�@      @                ��0=��?      @                M�nm2�     �m@                ��(��&�      .@�E�2	�?x}��Rs"@              �?��|��a@e��f��@        [9���?FB[Υx�?�p���@        J�=���?�;��)��?�$�A���?        f�"Qj�?                        ��ݮ��?     �C@M�'~�%@        ��E�Ը?�-��X@�X���?        .�u�y�?                @U2�s?�     �e@                9x�:@      .@                @U2�s?�     �e@                9x�:@      .@                ����G@      @                ��ve&�      5@                �%� ��'@      :@                ���<*@     �K@��6@�?�Ք�3�@              �?:@0G���?t��$�"@        �>�%C��?�x@�@�E��i@        �u�y��?      @��,5	[@        �������?     @A@F$��|@��P͚h��#Qj�a�?                �]O;@     @S@                ]���Kb��      @�G�z4Q@+��@        ��).��?      #@��+K��@r��S��?�Y@�H��?                E*����?      @                ���Џ�2�      <@      @^0�E���?        ��6�S\�?      )@                XG��).�?                &*�}�f6@      Y@                X-w���      B@                z;&����?      @                �	�0�     �A@                (��!R#�      3@                r�ޮ)�      4@��	ܺ��?�<�ǜ�@              �?�(�~�?�����@        ����o�?7�ُ��?a�H��@        E���Y@�?                �h$7�2�     �l@                ���+��      @                        ;ڼOqɀ?      !@�;"�a�	@        �۵r�3�?                8|�9�@      @                M���G&@     �M@                9d�(��      @                [U���+@     �K@��ʡ-@@5�+�H@              �?      @>��s��@        j�a�/�?��H�=�?�|��T@        �g�t�?��&����?                #Qj�a�?�G�z41@n?�=�?        C��6�S�?p_���?R?x�7C�?        5�0��?�!�uq��?�ү�@        ���o��?                S�u�l+�     @\@                �1��E�      @                ���@      @                �^/��3@     �a@                d�O��V7@      W@                L`n���?     �K@                ��0�+�      @                ��.�a�.�      9@ɫs���?�@���`@              �?^��K�?���C�=@        ��}�K��?\�C��@�|�7�@        �d����?                �S���(�     �l@                �pP����      @                �Fpt53@     �M@                p������      @�(\��:@^Ѡ�.=@              �?      �?'x�9�@        ާ�dֱ?+��^B@C�]\)u�?        �h�>��?                        ��ݮ��?�G�z41@��`8o�?        �/�Ʈ?                �5z N!@      F@                ��Tw�      m@                �5z N!@      F@                ��Tw�      m@                �*��      @                T�����      (@     �<@>�4��@              �?      @�����F@        �|�(5��?     �6@�t_\@        ��]+'�?���1ZG�?i�SY�@        ��Y@�H�?     �L@6�n�L~ @        �D���?     �=@�H^�|��?        �y��!�?      M@\-��N@        #Qj�a�?                q���[ �?      @                �yp)��      <@     �E@t���v@        �0���?      R@m�N��L�?        ��!XG�?                I_�xW@      5@                s��&���      @                K���]@      @                ���av�!@      (@                &AW�j}@      @                ��\0�r�?       @     �1@�E�jx@        ����, �?                        j�a�/�?      )@	}[��@        �f�"�?�G�`�9�?�wAn|�@        ������?                ��M@      5@                }���h*G�     �g@                Ҙ�Eb�      @                �����#@      0@     �>@��2W
@�F�7gXп�, _$J�?,e�X�@	Et4��@        ��o��Z�?                Gut��`5�     �U@                ge�rU�<�     �I@                Ƨ:s�@      G@                �Q�	G�      @N�St$�?\�l� @              �?��Q��2@%���k@        ��Rc�?V-��F@���%�@        �t�VN�?                �˄�B@      @                ��xw�9�     �b@                G>�_�g�      <@                a�
A@     �]@���~�z�?�g�i@              �?��,`w�?��6��g@        ��:��?��C���?T3P��@        ���}�K�?      �?��d���@        p��Z9��?�Ws�`N�?v�
fa,�?        )5�0ȷ?                C �	�)@      9@                ��@     @R@                        �k�g�{?      '@���L@        ��D��?                ���}���      "@                ��l��"�      3@                ���}���      "@                ��l��"�      3@                ����2�     �]@                (9����@      J@�[Z�{�?��^l�@              �?      @���}q@        �g�t��?'�o|��?
b���k@        >��E��?                        �k�g�{?     �V@k�!\���?        ���}�K�?                        �"Qj�a�?�A�La�?�
:{M@        ��Y@�H�?                ��?�?@      @                dԛf!4@      f@                ��	m�8�     �[@                .��ڌ�?      @                ��	m�8�     �[@                .��ڌ�?      @      @@��A�ʡ@        ������?���Du�?W׊�p@        �ݮ��?     �2@D��ym�?        �Y@�H��?     �G@�B.*"�?        �/�Ʈ?��C��G@�oW&@        j�a�/�?-���w?@k���R@        q�����?                �<��?@       @                �^/M˕ʿ      <@                >t���
�      &@                �%� ��      @                k���s8@      @                b�f�?      @                �Ut�0��      @                z����
4@     �[@������?�tI��@              �?(�o|�Y�?�t�
�#@        Qj�a��?���B���?���}�@        ��	��7�?                K�67T5�     �b@                �8g��       @      "@���!�@        &C��6�?���Y@�l��N@        �g�t�?                �4�{	:�?      @                rЩ�b�)@      *@                �����     �M@                H�u	�(@      P@fffff�G@cL�Y��@              �?�����l3@�L *e�	@        �`mާ�?��v��rH@��ƅ�@        �Oq���?                ��J�|@      @                X��(�9�      [@JF��@                ;ڼOqɠ?bX9��O@}j��H�?        �u�y��?                �4�A/#&@     �d@                ���	�@      5@                ��{Z�     �U@                |�����-@     �W@      )@%���@              �?      @�E�;@        J�=���?     �;@�qo@        l�g��?fffff�J@�jːU@        �g�t��?z�G�rG@ 6���}@zT�:;��Z@�H��?���y���?5:�č�?        �"Qj�a�?     `R@qQc{�E @        <�ߠ۵�?                �	s�R@      @                ��[e @      @                ���!*@      S@                �j-�@      &@                ,�ts��      ,@                �l��ƅ@      @                ���|ɉ7�      V@                �B��"@     �W@�o%;��?ĩ7ް! @              �?������?��Q%�O@        0��f�?��Q�h�?��
�R@        �۵r�3�?�O��n�?�y6�a�?        �(5�0�?     �F@��}@        ��ݮ�?                ��*� @      "@                �l���0@     @_@                ��u�(�4�     �`@                ��_!�      3@                *G"vq�      @                r��cm @       @     �9@i�l�E@              �?      @��/)$@        *.�u��?     @C@ %{�� @        ������?      +@;�e^��?        ������?      +@q�E���?        �����?      Q@���T]
@        ;ڼOq��?     �L@�ҭx90@        �6�S\2�?                ��s��@      @                f��ԨJ�?      @                 �f���      G@                L�'C}�;�     �]@     �:@o���M��?        �}�K�`�?                        ;ڼOqɐ?     @J@f����	@        �g�t��?�� v���?����?        [9���?                D���Y¿      @                ��9�.@      4@                D���Y¿      @                ��9�.@      4@                1 ����?      6@                ށ�㌔�      @                P0�Q@       @                V�A�#@     �L@     @B@��\�#@              �?      @w��ms@        ������?��C�l�M@��ڇ��@        ��!XG�?                z�!�g@      "@                � l�^k#�     0p@\*����?���f�@        �0���?(\���Q@��&��?        Sc��|�?                ��L6*@      $@                ��;L`�@       @                ��r0��      @                -�Ym@      "@     �Y@�E�]�@              �?�I�5�/�?�1�L��@        [9���?     �^@]h����?        )5�0ȷ?      K@��Q+?}@        ��o���?     �2@��+�K@        �6�S\2�?                �o ʋ�#@      ,@                LЦ�N�@      1@     �@@v;���@tk�P\���h�>��?      O@���+�4@        #Qj�a�?                        �k�g��?     �d@�N�t<@        1��R�?                �AJs��      @                ��� �1@     �R@      -@P�yF�B�?        �=��E�?                        ;ڼOqɐ?                �5*�@      @                gQ�9�1@     �P@                �5*�@      @                gQ�9�1@     �P@                ���>&�$�      T@                
��1�      @@                ~ؕB@      4@                Ε����     �M@      +@'q6!�@              �?J��&�?�Bh�@        [9���?     �D@S��f�@        ���Y@��?                Q��T4�     @P@                z%���@      (@     �A@�^Z8�@        �k�g��?     �<@jib��~@        ��Rc�?                �c�/@      d@                �<v�ɺ�      3@                �H�Gi�@      ;@                �.uy .@      0@     �8@P�JK�1@              �?      @�o��@        ;ڼOq��?     �9@��z���@        �K�`m�?                        �k�g��?     `\@8���l�@        �D���Y�?q $���?,���@        #Qj�a�?     �N@����>Y @        f�"Qj�?                LE'��y @      &@                �|���@     �`@                �I0��@�      b@                (�s��@      @                3���r@      @                �Mk�?      @                Ц+O#@     @`@                j^м�      @      )@�@BR]�@              �? �rh�]G@��)��@        J�=���?     �>@����@        l�g��?      @TY*A+�@        ���}�K�?l����J@:�^Fq
@        �H�{��?                !-��9@      W@                �XXr�7�      @                y�(�F)�?      5@                �"jc�L>�     �Q@                ���Q�2"@      ;@                ��;����      U@V-��F@�����"@              �?     �2@JlY���@        �	��7��?     �1@���Q@        {���?                        )5�0ȗ?�G�z41@��iv��@        x��A�k�?      G@�)n@        �}�K�`�?����B��?^,���g@        +'<�ߠ�?                �Z%(S�"@      (@                T=s ٙ<@     �g@                �Ry���      @                �k��<S2�      W@                �≬`���      @                ��=n&@      "@                 ��3^-��      T@                �5���=@      [@Ȱ�72��?��0� @              �?l�]h�S�?U�L��@        Nx��A��?�G�zN<@&X-H@        c��|��?     �N@k�=���@        �h�>�%�?vۅ�:��?�no&v�?        j�a�/�?                �L��
@      @                .�c2�Y4@     @\@      @BV�- �@        �Y@�H��?                        j�a�/�?                r�'�      @                )�p�f�      @                �P�Е @      @                �^����9�     �d@                �P�Е @      @                �^����9�     �d@     �V@���e�"@              �?O���|��?�r\�s@        ��!XG�?     �4@�>��V�@        �u�y���?                $�X�A�     �d@                -`aA#G&@     �U@     �\@�S����?        j�a�/�?      7@�icyH� @        �7�v���?                *�N@      @                �ǢE�@      @                ۃ�Tj���      @                ng�[&@      B@     �A@�3����"@              �?      @�~̇�7@        �۵r��?     �5@�!�%�'@        �|�(5��?                �#3��@      $@                ~�$�S:�     0p@                �hD^��?      .@                x��Gd,@      .@2���#�?��h @              �?�)W��?�� �B @        C��6�S�?r�Z|
 @�eŷvg@        z��!X�?                扶��n<�      g@                � !D��"�      3@                {�4�V"@      4@                d��%ʯ@      S@     �Y@�[��.@              �?      @�mH�}�?        [9���?     �^@��5آ� @        )5�0ȷ?                B�*Z��@      >@                �u��&�     �n@\*����?,u����?        ��ݮ��?     �c@0"�����?        �k�g��?                V��U(�@      @                ŗA�8�@      @                ���v��?      &@                tx���@      @     �<@�j���@              �?     �9@,�¢�1@        �|�(5��?     �F@���ҔA@        ��]+'�?                �Z����?     �h@                J�w9$�      5@                %��=S�     �@@                �3��7@      G@     �2@3q�,�@              �?      !@��k iN�?        8�v����?     �4@t���@@        @�H�{�?                g3��5�     @[@                ������     �d@HĔH�W�?D<,��v�?        �"Qj�a�?     �4@�4���?        �u�y��?                �áI@      @                "?v��� @      @                ��͊�q@      $@                ���f��      @      @
y�@              �?�=�>tA�?:���@        �����?     �8@��5f@        ?�%C���?                Ӳ�Xd�@      @                ���?      @      <@�8�,��@        �>�%C��?     �N@��*��
@        �K�`m�?     �0@�204$N@        �����?     �1@�~��:��?        �K�`m�?                (�i$$4@     �a@                J�hR�q�      @     �<@Y,1>��@        ��|�(5�?     �8@�&R�8��?        o��	���?                �iۥ�n@      3@                ���!|��      *@     �9@��t�
@        >��E��?Q�|a��?                XG��).�?                z,خ|5�      E@                ���s�� �      0@(��y�?p��+8;@        T\2�h�?                        ��ݮ��?                7`aA��@     �E@                y8�s�?      @      !@9���K@        �k�g��?�St$��?`�M\c�?        ��ݮ�?                �������      ?@                ��^�<@      (@                "�9 @      @                ' /��s �      <@                �*�g;�@      @                �OcUE�@      "@�7��@�.���[@              �?^�}t��@�&v_�@        i�>�%C�?     �8@j�$k��?        \2�h��?                pd��j�&�     �j@                ���.:�      $@                ,�8�4@     �Q@                |K�@��      @     �C@�K %� @              �?     �W@��L�@        G��).�?��MbA@jkh��@        �!XG��?                I��+7�     �k@                N<�`bB$@      :@�ׁsF @                �Y@�H��?R���AD@���RA�?        ��Y@�H�?                i��p�B2@      G@                ���r�\ @      @                �=���,��      @                �~Z�+@     �D@�-�����?�m�Zz�@              �?������?H3��2�@        0��f�?���[f�?�"���@        �۵r�3�?     �>@£ �M@        ݮ����?�A�La�?p�45�1�?        �����?*������?ހ�"��?        ������?�[Ɏ�@�?�V� @        �{���?                �{Sf��?      @                ��Y�9Y@      @                �޺�j� �      @                ���g0@      `@      0@��gS��@        ��d���?      J@��K�1@        j�a�/�?                Jo��8�      &@                ��b��%�      @
.V�`��?�wA"�A�?        ��ݮ�?��g\8��?}P�~�@        l�g��?e�,�i��?�Z^#8�?        �7�v���?      -@                XG��).�?                ���b��      3@                �YS��%�      0@                �=$[��#�      0@                ���!�      3@                >�T�4g�      @                �	?,���      @
ףp=*E@�
��O�@        <�ߠ۵�?     �6@%�g�"�@        �"Qj�a�?                r%a+��      9@                I��H�I&@      M@                𹸨R3�?      @                 �����@      @���e%�?og��C�@              �?�T�t<f�?(\���	@        �۵r�3�?,e�X�@�V_�B�?        �H�{��?c�tv2x�?,e��@        amާ��?                        �/�Ǝ?                ���x5@     �Z@                �!|��L�      @                ��]i�}:�      f@                �?W0pU@      @                ��]i�}:�      f@                �?W0pU@      @z�G��?0"��E @              �?�����	U@n�K��@        �d����?^�/��?uHk��� @        �6�S\2�?                ��4��     �d@                ����Tg0�     �A@                ���M�#@      3@                �?�Z��&@     �S@��� #@dQ����@              �?�0���?�Is��@        Qj�a��?      B@��V�y�@        �k�g��?�E�2	�?�ѡ�`�!@        ݮ���?�������?�����@        )5�0��?                vQ��l��      @                u���l���      @                ��XG-;�     �e@                3�, 1@      M@                �c���5'@      6@                v����s@     �B@      @��@ 7@              �?z�G�P@�����?        �g�t��?��� #@�ͤ�@�@        ��|�(�?                ����%�      3@                ���s��      @w;S���?�;w�t�@        amާ��?      %@��V�y�@        �k�g��?(�rE�?E!K���?        L�`m��? �J�R�?h��R�}�?        T\2�h�?                        �"Qj�av?                        ;ڼOqɀ?;S��?*N��3@        �H�{��?���`�?��
��@        j�a�/�?                Z_�d�@      @                +��v�t&@     �E@                Z_�d�@      @                +��v�t&@     �E@                Z_�d�@      @                +��v�t&@     �E@`q8��?d���_@        ��|�(�?                        �k�g��?body�?����S�?        ��ݮ�?      %@��#MB��?        �}�K�`�?                �ƾx�      "@                "�KFy��      @                A��%@      @                �@Ƣ
�?       @      @w��@        0��f�?V���n��?;���q@V�æf�?�S\2��?                Ѫ��<�(�     �R@                u߭}�5@     �]@                ��z@      @                �p�m�0�     �Q@                        �"Qj�a�?�f����?���]'@        ��	��7�?                �曡<�@      @                �3�
]�/@     �\@                (��N��      <@                j�IoO�3@     �U@��yS���?�nѽ�@              �?�ܵ�|��?D(��@        �Z9���?��Y����?M@�Ob@        �Rc���?�-�l���?�l{��@        UUUUUU�?�����?                �Y@�H��?                �r��"@      @                ��"�$�0@     �e@                �l�j(>�     �[@                派��
@      @                ϱMl,7�      [@                �#!�      @      -@7����Z@              �?      5@��6�!�@        �S\2��?     @B@?-���@        ���}��?                H<q��6�      N@                MJ�(�@      L@     �9@&D���$@        E���Y@�?     �D@3��V(�@        ��D��?                 �!�\;@      D@                -��xI�@     @W@                L]�&HE!�      3@                ��+ ��?      ?@�c*���?߲�+�N@              �?p=
ף�U@;����X@        8�v����?q=
ף0�?#�j�4N�?        �/���?                E���r�-�      h@                &�@�q�      @                ����>�@      .@                Ǔi!@      U@     �@@��+�@              �?      @�إ�h@        T\2�h�?     �E@�N����?        ��6�S\�?N֨�h4�?�X��[�@        �k�g��?��6@�?�*�~�@        ݮ����?                "L�o~�%@      5@                �7����?      *@                ��P
�7�      $@                �D��.m(@      >@      I@�fD�;@        ��f�?      !@�)b4�4�?        +'<�ߠ�?                T�g��h:�     �S@                 �oyA�?      T@                �4�c��      @                ��!�=+@      P@��\���?O�[@              �?7���a�??�@        �Rc��?GɫsH�?[׼�Ha@        �۵r�3�?R'�����?�����@        t�VNx�?�D���?D���@        ާ�dֱ?'"�*�?                )5�0ȗ?Cs�FZ
@ {I���?        ���:�?                ��,z�@      (@                ���JMM)@      M@                i����-@      N@                ��|L��      @                ��t7�� �     `f@                ,��oiS@      8@|�/L�J�?�K�`g�?        ������?M֨�(�?�XOĐ�?        XG��).�?                ���y���      @                ǫ-�y��      @                �C��E�      @                _�,"@      &@��jHܣ�?>^�a�"@              �?      @$�4�@        �h�>��?��?��?E��4=�?        �).�u�?     �E@�{Ƶ"q@        ��ݮ��?     �X@i :f�@        {���?                ��L�M(@      @                [�~m65@     �W@                �C�*u!@      @                x��.��      @                ��n<�YC�     �d@                9R._��@      4@     �K@�Y��<g@              �?/Q�5�U�? ��sb@        �>�%C��?�#EdX�?�6��5�@        �u�y��?                N9Nu�     �T@                y�I�q@@      `@     �Z@bz� ��?        ��Y@�H�?!����=�?:��e�?        �|�(5��?                	��H�o"�     �@@                �z�� &�      0@                G+���@      @                ����S�@     �A@     �0@[|nz�@              �?      @��CEEp@        p��Z9��?     �X@�jg���?        �D����?      *@k�d�E�?        ������?���ت�?�o�a@        WNx��A�?      -@X�#@        �7�v���?                        �}�K�`�?                �E|јw@      @                P���DE̿      @j�t��?�*L"�@        .�u�y�?t{Ic�
@#�ۜہ�?        �ݮ��?      6@��z�t�?        XG��).�?d�CԷ�?                XG��).�?                ��n;7��?      @                ��p7%�?      @                W�ɵ&(�      5@                M4��L'�      @                ɟ�&ϰ$�      5@                N�ým��      @     �C@s��@��?        v�y���?     �B@�x���g@        t�VNx��?                ��Xb52@      V@                ��" 2�     @d@                �X��#@     �Q@                �� @      2@     �;@@s��4@        �"Qj�a�?     �C@ێvn��?        �0���?     �?@!+��@        �/�ƾ?�VC���?/�y�"@        �}�K�`�?                K�l$���      @                Ί��"�      B@                ���,@      <@                �wG���@      &@��h oA�?Ѝ=��j@9�߳8����D��?�k�)�@����;��?        ��L�n�?                -+�ȃ1�      I@                x��FB�      @                 �+�@      *@                ��č-�@      .@\���(�H@��)#�@              �?�_{f	�?j�,�)@        �).�u�?     �U@m�W��@        �h�>��?                DKS���:�     �W@                �\&��A@      @     �B@t&4i�f@        *.�u��?�p=
�CJ@�Щ4d @        i�>�%C�?�G�zNL@���{@        �|�(5��?)\����V@d����@        ��o���?                ��k@      @                '���#@      ?@                Oſ� �@      @                +п�Ż@      @@                �O�~0�     �S@                А�:��@     �H@      -@a���@              �?�x�&1��?�s)cd�@        �S\2��?     �4@�+D��(@        ���}��?      @���R�@        �=��E�?[rP�@�b 1��?        �Y@�H��?                E]m� <@     �]@                �:frA�?      R@                Wq���z@      $@                2��v�V<�     @R@                �.�@      @                ��pu@      2@     `Z@Z{���@              �?     �5@��D�i��?        4��]+�?      2@�I˸��?        �Y@�H��?      %@�)��Nv�?        �h�>��?��H�}�?F��@        ��Y@�H�?                �Qf���?      @                [�f�@      @                ^	�5�@      *@                �Q�>y'�      U@     @M@vs(���@        �}�K�`�?F���j�?����@        p��Z9��?                ���Ա/@     �Q@                @W�P)@      @                ���J�
*�     �I@                ���ު�#@     @Q@     �g@�����I@              �?     �K@��En�9�?        �!XG��?                        XG��).�?     �A@����i@        ��|�(�?     `R@�0���"�?        ��ݮ��?                ��,E['�     @q@                W�:V@      3@���ڧ��?E���`u@        ��d���?     @B@�c6�q@        ��o��Z�?                �a��p�@      "@                `��zW���      $@                ����T�*�     @_@                
�}k<..@      U@�yS�
#�?�;3h @        �/�Ʈ?     �Q@�v���u@        ��D��?                V>�e�T�      *@                �Ĵ�g��      @                �>�
s��     �F@                �⬰��@      @���ڧ��?�i��o@              �?     �:@�t��I"@        f�"Qj�?��<�!� @g���aL@        4��]+�?                ���Z=�      f@                :�\�'!@      &@                �.&O*@      ;@                �3�π>@      U@     �T@^�4y��@              �?     �S@;p_5��?        M�n���?     �4@��gsn@        ��E���?                �E�C��*�     �l@                ���ؠg�      "@-C��6�?                �"Qj�a�?     �2@���jZ�@        mާ�d�?                �U�͎-@     �A@                ��j�jJ@      8@                ���Q,�      0@                -��3q-@     �B@     �<@��r��>@              �?�vö��?��y�=]@        +'<�ߠ�?     �1@ <��r�@        ���Y@��?     �;@i�EQܘ@        ��o��Z�?     pe@}O�u��@        q�����?                p+f�?Q�     @Q@                2�-S6@      O@      ,@�v���?        Z@�H��?      '@�k2�@�*�}��׿�!XG��?                ts۔*@      K@                �:
����      @                �D����	�      @                =�����@      I@                ��L0�e�      *@                ����R�7�     �D@      G@���{շ@              �?p_���?���i@        s�3���?     �4@eX��@        �f�"�?       @�3M���?        t�VNx�?     �2@p��z��?        [9���?      M@�����-@        >��E��?     �D@Z~��ua@        ~�K�`�?                ����#�      4@                Y2&�/�     �U@                k��[��      @                �zV?�#@      A@                h�L,S�?      @                �Q��+@      2@                R�k��     �[@                +ާ��'@      6@��jL�?d}��@              �?     �R@��O��@        >��E��?T�t<f��?����@$@        �g�t��?     �1@̣0��@        9����?     �2@"s$��r!@        �n��	��?ܺ��:��?^��C�?        '<�ߠ��?                        �k�g��?                ��+U;+,@      A@                �����#@     �R@                ��+U;+,@      A@                �����#@     �R@                9����>�     @T@                ���Cy�@      M@                P��hP�      6@                ��?��-@      :@      !@7�%|@              �?��+H��?%�����?        j�a�/�?
ףp=zF@��3=�@        9����?                D�$i%�@      @                `"<lN @      @��<�!� @g����@        ��A�k��?     �2@=
�^�@        f�"Qj�?     �:@����@        �u�y��?      ,@���cV��?        j�a�/�?     @K@h�)@        ��, _$�?
ףp=�I@���P4@        �}�K�`�?-��阮=@�z�?        Sc��|�?                        j�a�/�?                �;8�-�      @                {��i��      @                 ��%f#�      3@                �ElS��!�      L@                 ��%f#�      3@                �ElS��!�      L@n���9H@������@�$N����?t�VNx�?ޓ��Z� @'�y���@        �}�K�`�?                �%}�cL@      $@                �M/+0q&�     �Q@                ��3�R@       @                #�y�0@     �W@ �rh�MN@<�m��?        �/�ƞ?2ı.nc@sҨ��?        �k�g��?                �~��EM�      @                �������      @                ��"����?      @                �|����?      @     �0@B}~ш�@              �?     �9@w9�L�@        <�ߠ۵�?     �5@��Yƴ��?        ��|�(�?     �:@��8��@        _$J�=��?�#�G[�?	��\� @        �:ڼO�?                ⸥ܚ�0@      D@                hYǹ���?      *@                bWEj��@     �T@                F�?j#@      @��6 �?��֤�@        l�g��?!�rh��D@(�D]�@        [9���?                2!F�/A8�     �T@                �����R"�      &@                
��)z@�      @                C�A<�%@      N@2��*��?�Gq@              �?4�Op���?,�5��)@        c��|��?     @N@��*Ѳ^@        s�3���?     �D@0�{
�1@        ��ݮ�?     @D@i�	�@        �����?                �[�Ծ\0@     �K@                ��Ӑ��      (@fffffT@���D�@        XG��).�?�/�$�Q@ ���O@        $J�=��?                ����U)�      1@                p��N���?      @                .�T:�B�     �b@                fN�cJ@      (@      >@��"�@        �}�K�`�?     �T@E�����?        �Y@�H��?     �K@�[;a� @        �u�y��?      C@�-���@        &C��6�?                ��
_���      @                �Kzͺ�      @                ��h��8�       @                �J�V��?       @                
;� �/@      .@                �;��?      $@     �5@&T��I@              �?      9@"ǅ�1@        ��A�k��?&1�Z�?+��3�I@        ��E�Ը?      )@-LU77��?        )5�0ȷ?      +@Ɠ��<r@        �"Qj��?      1@6L��7�?        ��ݮ��?                        ������?                �B0 Y@      @                ���Eg!@      8@     @`@arTC���?        �D���Y�?      %@���M$@        �VNx���?                RV�6�0�     @R@                c��Q� @      @     �1@                )5�0ȗ?     �0@A�R� @        ��f�?                &r�߿      @                �ċ�Wr$�      *@                &r�߿      @                �ċ�Wr$�      *@                a������      @                7{}�6��      $@                �΄RK�1@     �K@                d���"@     �[@���[�?�n6M�|@              �?N֨�h4�?jQ.��@        B�k�g�?�?��"�@�qD}{L@        }�(5�0�?                �F:/"�     �d@                ���6��      $@                �g+��0@      I@                ��	l�-@      R@     �8@PV8WA@              �?     �1@���	s]@        ;ڼOq��?     �9@ciJ��@        �K�`m�?                B"�m
�     @Z@                q-${-�0�      J@     �2@�˰F� @        #Qj�a�?     @L@5�K���?        f�"Qj�?                NCYF��@      @                �F��_ @       @                P��F� @     @]@                	�u"@      (@����^u@H���ɥ@              �?��&��O�?�%k��/@        ݮ����?b���i@\�"����?        F����,�?�2��bb @5��z�e@        �K�`m�? o���?��Թ�@        )5�0ȧ?                �&xxj	@      @                k��%@     �R@H��Q,7�?k���[@        J�=���?                        �/�Ǝ?                        �"Qj�av?֭���w�?�Zeb+�?        ������?                Y�IQ\,@      @                ��3lG/�?      $@                �*��&Կ      @                :"�'2�?      @                OA�H~A�     `h@                !�!+�v@      @                OA�H~A�     `h@                !�!+�v@      @      +@z�,l @              �?     �4@�h�a�@        ��ݮ��?      4@���/ �?        ��E���?                Z������?     �c@                I�D-��(�      <@                ������1@      L@                i� �}@      M@     �8@s#σY@              �?      -@��&���?        q�����?�j��� �?rq�շ=@        ;ڼOq��?�ʄ_�g @���%@        �S\2��?     @A@�oj@        �>�%C��?     �5@���h�u@        �ݮ��?�bE��@����e�?        �0���?�'I�L��?                ;ڼOqɐ?     �:@��H(��?        ��ݮ�?                ���.�      @                4�*��U@      6@                �6"- o�      @                ��O��@      4@                |ݩ�� @      @                F��L�/'@      "@�-�����?����s@�P��D����ߠ۵r�?���խ�@5��1���?        p��Z9�?�=�$@��?�Z.��@        B�k�g�?     �F@���H�F@        �f�"�?                �p!�� �     �N@                �5��'(�      6@                8�����@      @                d����r@      ;@                >�
y�$�      W@                l/LG�V!@      <@                �_/��%@      (@                ǦS��       @
ףp=zF@�ֳ;3@              �?     �0@L���X�@        �/���?���Mb�F@v[�4Z�?        8�v����?     �F@�wm�`�@        �۵r��?      6@�Ѹ��q�?        �u�y��?                �q����@      @                uRz,�0@     `g@�=���d�?����٤@&݈��ɿ��Rc�?                        �"Qj�a�?                ���`�@      @                83F)��?      @     @Y@��ڹ�M@        j�a�/�?                        �k�g��?                h��8J:�      V@                �?t*��      @                ]l�[<�     �T@                �r�� @      @                ]l�[<�     �T@                �r�� @      @     �Y@S:�ۚ<!@              �?     �?@����0�@        [9���?     �[@�4~P��?        )5�0ȷ?      @+�!�@        f�"Qj�?9�ֿ@                ��ݮ��?                U~��v�@      @                
yޗ��&@      :@      (@��UO--�?        ������?     �8@்w@        Z@�H��?                �c�/V`
�     p@                ��L���      @                W��o�U@      @                j�Lcj@      $@     �9@�xxf!@        �g�t�?     �=@��x�@        �����?                ����h�:�      W@                �@�0�@     �B@                �44�"@      B@                @
1���     �T@      �?�m;���@              �?      8@�V�~���?        #Qj�a�?     �8@W`p��/
@        �Z9���?                �����i@      @                �'SRH@      @                � �C�=�     �d@                U|.@      `@�8�ߡ��?gT��@              �?      /@�����@        b�/��?��67�'�?��8y��?        <�ߠ۵�?                XC9��)@     @U@                G��b6�8�     @`@                �rU�%@      7@                �[ߊ�{ @     �N@��bE��??���@              �?l�`q83�?C�i�H@        �"Qj��?&�lscz@�ܾk3 �?        �t�VN�?�0�����?����=	@        ���Y@��?      @)��,:/@        �u�y��?                %/웢M@      4@                �ILr@     �B@�=yX�5�?9��h�,@        t�VNx�?���7�v�?n��|Z0�?        j�a�/�?                        �k�g�{?                        �/�ƞ?                ��>�0e�?      @                �[fVp��      @                ��>�0e�?      @                �[fVp��      @                z��wG�A�     �i@                s�f&��      @                j߀dO[@      @                �n��k��?      .@      @���( @              �?      @G�N_;K@        +'<�ߠ�?�G�z�0@�Hg�3.@        {���?                t���a"@      @                ��7b� @      4@                ���4x@      @                 5蔐��     �p@     �1@��8>l!@              �?      @J�o�@        ��o��Z�?     @Z@K��y�@        1��R�?                <򧵳J�?      @                F�k,�:�     �Y@     �J@ؐF��w@        {��D�?      :@P��կa@        ����o�?                �v���F5@     �a@                �_��Q!�      @@                =�9�',"@      "@                �������?      &@      @A�"SMA@              �?      @�����h�?        ;ڼOqɐ?     @@@ꢓ�T�@        .�u�y�?                8�o�6
�      @                �X�4��      @     �2@	�F�[�?        ���, _�?z�G�rG@��I�� @        �, _$J�?                ������?      =@                dS/Eo0@     �J@                %R�&�4�     �P@                �Z��@     �a@j�t�F@*_�f�@              �?     @D@��V�D@        ������?ףp=
L@���@        ��).��?      '@-c��Gs@        G��).�?��Q�>I@u�*�c5@        �����?                �E��{�/@     �M@                d������     �`@                <7�}>n�?      (@                ��5���?�     �S@                �	��D��      "@                vV(_��@      "@     �6@��]�W@              �?     �5@�|�+BN�?        �%C��6�?     @B@�����@        mާ�d�?                �?|)�     �_@                ���F~��      "@                y�OM�P9@      [@                ,��B\f�      L@R���F@�\1�M@              �?`��"ۉB@�4��-�@        �7�v���?�K7�A G@f�1��U@        �D���?                ��"�9��     �F@                bޕ{�&�      :@     �J@�*��q�
@        j�a�/�?+�R@ �� �o@        ����, �?                z6`��_@      @                V�(�M�?      @                ��8���     �Y@                ���+�4@      ]@     �X@�LR@              �?     �W@s@�{��?        f�"Qj�?      &@y�k�@5@        ��7�v��?                �A����5�     �p@                ܙ]
��      @                BX�)�      @                Jk�C!�+@      9@q�Ws� �?���x�e@              �?     �<@��`R@        ��Rc�?����}�?��4/��@        p��Z9��?���,N�?��F�?        e���}�?                        j�a�/�?                �bK�֜@      "@                �1A�%@     @`@                9#�57�      b@                'z���G�      &@                9#�57�      b@                'z���G�      &@� �����?��1Pϕ"@              �?��F��?���PB�@        j�a�/�?���8�?]��n@        WNx��A�?��e���?�8b��Q@        �o��Z9�?      3@�/Vפ�?        �/�ƞ?�׻?�?W!�J�M�?        �u�y��?�Z|
�q�?&L3��w�?        �0���?                ����-3(@      $@                �5���?      @                �Y3�xG��      @                ˙>@�@      ?@      #@8�c�R�@        &C��6��?�<I�f�?8en"ϣ�?        ��|�(�?                ����v��      @                է�Z���      @                0�LnL(@      $@                � �IA�     @f@                rt���@      @                f�[��"@      I@     @A@=��@ �@              �?     �>@	�mx��@        �D���?                        ��ݮ��?                ��y�0�3@     r@                Sf��g�      @                ��y�0�3@     r@                Sf��g�      @     �Y@`*x8�@              �?     �3@�k�y��@        [9���?     �^@��c��?        )5�0ȷ?                �/6��}/@     �c@                q���-�     @]@                ~��ICK @      &@                �?-[��@      ,@Է����?ᤕ�x@              �?      @�����@        l�g��?Ͻ��?߈��vi@        J�=���?                        �/�Ǝ?      C@T�'YG�@ЛY��ꉿ�h�>�%�?                O�6\=@      @                �����@     `i@                O�6\=@      @                �����@     `i@                cǪTry>�     �S@                ;��hi@      $@     `b@% ��v@              �?      I@��c�`U@        �%C��6�?     �5@�PJCcR�?        XG��).�?��n @�$� &@        mާ�d�?      /@�5ʦ�@        Pq����?                x�`Z�?      @                ��=EG�@      @                �Gl��� �     �a@                bQ�Q�r�      @                �ɹ��@      @                "i��@     �a@     �2@��^"�J@              �?     �0@{\��\�@        z��!X�?     �H@OZ����@        �:ڼO�?                v`Z�{8�?      e@                �9[���*@     �M@                ^�YnH5�      O@                (X�5��@      "@      +@�8��Q@              �?      �?D�LH�	@        ��ݮ��?     �4@/�X滆�?        ��E���?                        �"Qj�a�?     �0@��̏(@        �]+'<�?                ̊^Q�*@     �J@                N�e�#��?     �L@                ̊^Q�*@     �J@                N�e�#��?     �L@      !@q�����?        WNx��A�?      )@�ILTD@        �K�`m�?                l�W�B��      @                d-64՞�?     �[@                !���F�7�     �K@                <Vb��$�?      1@Ǻ����?� ^~�n@              �?     �V@>6���@        @�H�{�?���+�?<b���t�?        �ݮ��?     �1@]�p�O�@        2�h�>�?      F@_r���@        p��Z9�?                t��� @      @                l�����(@     �N@�%P��?=���g�?�L�v�ڢ�ݮ���?       @�I��^~@        ^+'<���?                ��'j)@      5@                ��&�b"�      ,@                $��7�;�      ]@                �-�� t�      (@                ��t����      @                ��P�~#@     �O@��MbH@��Y��@              �?���S�E@N����@        �:ڼOq�?NbX9�U@��v�LD�?        ��!XG�?     @Z@Y���V% @        �n��	��?VH�I���?U2Md�?        �0���?                ����*�5@     �a@                ��[d�      B@      K@�_���@        1��R�?                        )5�0ȗ?                �f�3W��      1@                *wk�      @                �ٸ�(/�     �L@                �e�]���?     �C@                �ٸ�(/�     �L@                �e�]���?     �C@      #@��t'@              �?     �9@A�M��@        +'<�ߠ�?     �1@4��
�?        {���?Qk�w�"�?v�_�צ�?        UUUUUU�?      @��<<|�@        XG��).�?                ��8��x�?      b@                �0�Ue�3@     �_@                ?��N�K�      0@                �<	J*��      @                *����M@      @                J�"����      @N�St$�?4?�x\@              �?$EdX���?�J&��?        ��Rc�?=
ףp�@@{�  A�@        �t�VN�?                ��9��](�      a@                <W����      @9��v��5@M҃�ͅ�?        ��ݮ�?�o��e1@'ǘ`�@        �d����?                �]Hm[��      @                v7LOu��       @                G�L�rN;@     �U@                �J�`�@     �L@
ףp=zF@��䷑@              �?     �=@�_
g�b@        �/���?V-��F@"5$��@        8�v����?      @Xt�?        UUUUUU�?�g?RD� @                XG��).�?                        XG��).�?      @I×Z#�@        {���?                F��E%��?      @                �Fp��4�     @X@                ݛ׻��.�      X@                ������      @                ݛ׻��.�      X@                ������      @}?5^�yH@�r��� �?        #Qj�a�?��x�@��?�.-uq@        �0���?                �~1����?      @                7�ATޖ#@      &@G�?��?���E�?        �=��E�?+��
[@<�R|� @        _$J�=��?                ˠ�Q�R�     �A@                �y"e*�     �C@                ګ@�f06@      X@                 8�.
�      @     @A@��Z�T�@              �?     �?@��%���@        �D���?                        ��ݮ��?���=���?F�h��Q@        4��]+�?                        ;ڼOqɐ?                �E�� �     0r@                &-��      @                {D��1�     @V@                YC�͛"@     @i@                {D��1�     @V@                YC�͛"@     @i@      #@�q��B�@              �?      @B"JΌ@        5�0��?      !@�a4���@        �g�t�?��(\��?@T��1$�@        v�y���?     �W@��$�@        �ݮ��?|~!<�?��r��?        ������?     �4@�[F��?g�R_4?��E���?                8Ӷ!�      3@                @~��@�?      @                ;P`�b�:@      `@                ���~> �      0@                �|�#�F@      1@                � �o��%�     �Q@                ���W�&�      B@                GC��(`�      @     �>@�5::^@              �?     �<@^z�ۜ�@        �Z9���?}iƢ�?Ԓ�R�V�?        #Qj�a�?      @�#Bv@        �D���?     �=@�Ց�=��?        �۵r�3�?                ��+����      @                �" Ժ��      @      +@8wxG��@        )5�0ȧ?     �8@Qw����@        ��|�(5�?                \ayۡ�@      @                �(4�-@     �P@      2@�$��2��?        �"Qj�a�?                        XG��).�?     �7@�T���@        ���}�K�?     @A@��DD@        �/���?`YiR
��?�J���b@�+g��.���VNx���?     �C@2	�@݁@        j�a�/�?     �7@17�p��@        �y��!�?     �7@�MN�@        l�g��?�'��?n�(z�9�?�tnC;ݿ�Y@�H��?:�}�k�@�˝�E�?        ާ�dֱ?     �0@�Z��r�?        ��Y@�H�?     �:@�(#��?        #Qj�a�?                q�;L�T@      @                ~\�7F@      @                "�,,��      @                ��`s�      @                =��|z9�      O@                פ7>��       @                ����N@      *@                j�Sg����      &@                ���x�� @      @                şw�T��      @                ���x�� @      @                şw�T��      @                ]�Su?-@     �E@                ��/-�9�      *@                O��^'�      @@                '�1V�@      @      �?i�����@              �?                        ;ڼOqɀ?     �7@'w�խ@        ��:ڼ�?                ��dk3@      @                �3v��     �r@�����?Tܸr�)@        �`mާ�?      @�լJ�@        T\2�h�?                ��+1&C;�     �W@                ���O��@      4@                �$��:�@      @                ���D�#@      f@      @2)\�$@              �?      @�k�L�C@        )5�0ȧ?      /@6�F�@        ���L��?                ���� T�?      @                ���F$�      .@      2@�5!�MH@        �/�ƞ?     @L@�i��Z��?        - _$J��?                        ;ڼOqɀ?      2@+�&'X��?        �"Qj�a�?                mŊ=��@      j@                F�}��!�     �N@                mŊ=��@      j@                F�}��!�     �N@                ��Ui��@      @                ��b���@      @     �<@�~�˞�@              �?     �6@#ӿ<:�@        mާ�d�?$]3�f��?�o ���@        �K�`m�?      @\�����@        L�`m��?     �6@����Ҿ�?        �S\2��?                t���Q� @      $@                �Kc�?/!@      L@                �f�z@      ,@                ��Tl>�     �X@                	�wnqS,@     @W@                ���yCI�      ;@     �Y@�ML�P�"@              �?      6@D9��B�?        [9���?     �[@�(p����?        )5�0ȷ?�(��?��QU�{@        �t�VN�?����?��?��F��@        \2�h��?                V:�s@      @                �;F~,(@      <@                ���"^�      F@                �f��E�#@      7@                r�mq=�      \@                b/�%��@      V@      -@bL7I @              �?      )@C��C^� @        ��o��Z�?�ek}�P�?6r�;�M@        ��D��?                �&�tJ]@      =@                ���\�7.@      <@     �Z@]c-@�@        p��Z9��?V0*���?ؿ��Z�@        ����, �?     �7@ ���v@        i�>�%C�?     �t@+$�����?        p��Z9�?                )u:"n@      @                �8�e4�@     �P@                h���!�4�     �Q@                032��c@      U@                �����%�      *@                ���
����      @     �5@Y�ǕX�!@              �?���QG@�"-;@        - _$J��?��d�z�?���8m7@        ��A�k��?                ϖʺ�%�     �R@                ��︦yC@      `@                E���+f6�     �P@                �4���q@      <@     @N@:z�%U@              �?      @��YG@        s�3���?      .@�qE-$U@        j�a�/�?                /j�Ok^@      @                $�o/�     @q@                        ��ݮ��?     @E@�T�<U@        .�u�y�?                aG�+`��      @                ی�D�)(@      1@     `R@���D�?        �k�g��?     �S@;��ͣp�?        Sc��|�?                b���Hd@      @                �
|��@      @                �������?      @                �o?�2H@      @      @b��j�@              �?     �1@?J��5@        �����?     �8@�v�W2) @        ?�%C���?                        �k�g��?R~R�S�?>�T���?        #Qj�a�?                W8/h}k0�      b@                Dw��g�@     �a@                W8/h}k0�      b@                Dw��g�@     �a@                U���@      @                �ȣ3�e@      @j�t�F@�Xr9�@              �?      -@�H[|��@        ������?��C�\K@��4hg�@        ��).��?      �?)`��)�@        v�y���?      @��"
@        ��!XG�?                >���ݐ1@      M@                �,`w�u@      b@                �0*1�� @      @                ^4���9�     �R@                �R�FE��      "@                &CB�@      "@     @A@����@              �?     �;@�W��'{@        �D���?                        ��ݮ��?      /@*��_T�?        ���o��?     �?@�����?        �ݮ��?                ���Oo@     �q@                K=���      *@                �A�G'@     �Q@                �BpB?��     �j@                ��brM(�      "@                 O��jJ�      @      %@���A�@              �?>
ףp�7@��H�8@        ��7�v��?     �4@�k���@        ��E���?                        ��ݮ��?���	���?M$N�N@        ���:�?                �1�A4@     @R@                0s�K�_Ϳ     �d@                �1�A4@     @R@                0s�K�_Ϳ     �d@���gV�?�\W�`��?��W-���<�ߠ۵�?�`��ü@�˩����?        �ݮ��?                ������0�     �C@                ���8T��      @                �4Yt�@      "@                ��4�$��      @     �I@j~F��@              �?{�G��Z@6TH���@        M�n���?     @L@��Խ[�@        ��E���?     �1@�qA+@        �|�(5��?�F=D�{�?                �Y@�H��?                2Xۚۉ'�      :@                l)���ſ     �B@                ��l���     �W@                ��c�,�@@     �`@                ;�B��@@     �h@                �R����?     �@@��jL�?��<��@              �?      U@Y��ar@        >��E��?���=���?�����?        �g�t��?                �3j���2�      f@                -����A*�      1@                �~�s�!@      8@                TlG��@     �T@      @��W��@              �?     �1@�!��<�?        ������?      3@��X��A@        z��!X�?                ���_�%@      @                J���8@      @     �=@`?��@        ��}�K��?�|~!�?���/� @        �����?      (@��'ڀ	@        �k�g��?�E���$F@��"��
@�"�ԡ�ӿ�r�3��?��Y����?�E��@        �E����?M֨���?�V^^�
@        f�"Q�?                �^�t1��      T@                ��W�]&�      "@      @��Rvg�@        ������?.�;1���?y��9�?        ��f�?                9�S��e@      "@                �G�{X��      "@n����D@��چ��@        &C��6�?�ʦ\! @J?
m��	@        #Qj�a�?                ��	G)!�      4@                .��_T�      @                t��6�� �      6@                �p�r��@      6@                8ւk�J��      @                ���%�$@       @                ���s(���      @                o�rI��7@     �Y@      @@�����@              �?      -@y����X�?        [9���?     �R@��.�@        ���Y@��?                �a:KG�@      @                ���P��*@      L@                ���j�2�      j@                �[�a@      >@      �?&��O@              �?                        ;ڼOqɀ?      >@���c�@        ��:ڼ�?                �Zm�@�@      @                ���D[?�     �r@���3K��?Z�j�@        �:ڼO�?      -@�8�6���?        �����?     @G@�:,@        �]+'<��?�� �B�?                �"Qj�a�?                w�!�Vy2@      e@                3������      G@                Oj���-�      J@                �=N?	�@      7@                �W�.@Z&�     �P@                �PD�� @       @&ǝ��z�?R�=��@              �?^����?p��L�@        ��	��7�?3��bbs�?Q��Ν@        ����, �?                mA�Y�.'@     �k@                �D�̫+@      @                3�����1�     �@@                ~_k=	@     �C@�x�S�?����U@              �?���S�e9@}�J�)K@        e���}�?H�`๷�?:D�?!�@        7�S\2�?43333�6@u�X@        ��ݮ�?�$���T@0G����?        �f�"�?                h�=ME@      @                �^�)@     �`@                t3���      $@                 ��ɭ@      @                �G����5�      `@                n&n��2 �      0@     �<@���>$g@              �?      @a�7�v�@        �|�(5��?      V@�p�9^H@        ��]+'�?                \��v�@      1@                �=m��l:�     `k@     �2@ �FA�"@        Z@�H��?                        ;ڼOqɀ?                ~��	�2@      A@                �,��{�      8@                ~��	�2@      A@                �,��{�      8@     �?@�M?Uچ@              �?      @����@        4��]+�?                        �Y@�H��?      )@>���>�?        ��7�v��?      P@�"�{��@        �}�K�`�?                ��ʼ#@      4@                lQf:�J @      q@                [+B��?       @                ���h�!@      (@�-�����? ,�C@        ������?V}��b?�?                XG��).�?                ����7%�     �a@                lё6@     �_@                �tWz|��     �e@                ���yZ,@     @W@�E���$F@�t�=@              �?����~��?d̻0�@        2�h�>�?�x�&1 K@�Ryz�#@        �}�K�`�?�.4�i$�?�c���b@        ��D��?��� ���?X�ƭ+O�?        ��7�v��?                hz�6�72@      K@                ���+�#@     �`@                &}�v�?'�     �T@                ��"�i@      *@                �7�H�y�      (@                A-.�LV�      @     @D@�����@              �?      @J���Q@        Z@�H��?     �C@��D;@        ��ݮ��?     �@@u�2\4;�?        ��6�S\�?      A@�B�5Ѕ@        �"Qj��?                L��W�*@     �D@                ��lH#@      &@                �/!?f8�      Q@                N��F\�?      (@������?D�b��@        mާ�d�?     �4@N��*3$@        ��E���?                �I��b�-�      B@                ��G��@      ,@                ��� hm,@      0@                � �£.@     @Y@�@��_��?e��
�@              �?      �?�3x;C@        ������?!����=�?�� �T@        mާ�d�?                        �k�g�{?     �3@ņ��d�?        �E�����?                ��6��y.@     �B@                �:�/�=@     @S@                ��6��y.@     �B@                �:�/�=@     @S@                g��K�'�     �e@                vɴ���      $@      @�Q���@              �?3�}ƅ�?���=�@        �����?5^�I:G@/��x]�@        ?�%C���?                �j�:�@      @                Ֆ��?B�?      @�Q��{A@a� ��@        UUUUUU�?     �9@�ɧ�@        �{���?                ;Ʝ��     �H@                � R�N�5�      I@                W��qQ,@     @d@                ��B��9&�      9@     �5@o ��@              �?      @�C۽���?        ��A�k��?��� � @1Cc�
@        ��E�Ը?                W�ܙ]Q@      @                � D�U2@     pp@                �m(��&�      4@                �s%�:�?      *@      /@`4x�l*@              �?      @��݂a_@        t�VNx�?     �D@\�㔙@        �E�����?                ��7Jw��?     �B@                &6P6�2�     @Q@     �B@�i?Bc@        �(5�0�?     �E@l�O'@        �u�y���?                �Q�3�Y@      b@                l�Q����       @                        ��ݮ��?     �G@#���@        ����o�?                7�X��@      @                ����'@     �B@                xx�X9�      @                Ȑ��#n,@      @@     �G@�%��@              �?     �<@c����@        l�g��?     �J@� 8]��?        )5�0��?D�+j�?��^��@        ����o�?�G�zN<@��8�84@        )5�0��?                ��o��!�      4@                }�sr�(�      W@      -@Ј$�n$�?        �]+'<�?�+jp�?���&�?        ��!XG�?                �u���      "@                �x՞��6@      Y@                �_^���?      @                K-�µl/�     �A@                �{<F��@      @                v<z��@     �@@     �0@0 TKĥ@              �?t���.�?E���9@        ��o��Z�?     �7@�16��$�?        �, _$J�?                Un+_��(�      R@                ~����l6@      X@                ���+�2�     �Z@                � �VW�&�      9@     �7@hg���@              �?      ^@Z�)2��@        �S\2��?      @��"@        ���}��?                ��02�      \@                +�<����      @      2@Y�.�@        ��E�Ը?      @�|�|]@        ����o�?      @'JѼ�?        ��Y@�H�?     �6@�sq{���?        �}�K�`�?                ��K�'�     �@@                �V�W�!@     �_@                0��L��?      @                ���%@       @                ����H��?      @                �Ʃ�i �      @V�`��?���^@              �?0�AC���?uȐp_�@        ~�K�`�?��n��� @O��5#,�?        �h�>��?�O��n��?���Gs@        ��f��?�H�����?�w��@        �f�"�?                ǁ���� @      4@                �~����@     @S@                ��`c�{-�     @e@                L��8�@      &@                Q����7&�      0@                h*w��z@      @��n���?�8��M@              �?���"��?9ޣԽ@        ��Rc�?����"�?U��K`
@        �t�VN�?��(\��?@G��s�@        9����?                        ;ڼOqɀ?                0=y�/@      @                �WC<�j(@     �b@R���1;@�tB�@        XG��).�?���S�S@�gq	�?        c��|��?                !�_�G@      ?@                O�d�=�     �[@                �� `\%�      3@                n��;�( @      (@                ����h"?�     �Y@                �-�B��?      "@     �Y@���p@              �?�(�'��?l�>�_@        [9���?     �2@E�"M @        )5�0ȷ?                E���;3�      c@                ��?�b�,@     �\@      #@b]�Y�@        .�u�y�?     �5@����?        #Qj�a�?                �D���.@      .@                0�r��      @                �����?      @                �n��J,��      @     �1@�,t@              �?���EB��?�rٙ$k@        ��o��Z�?     �I@x�����@        1��R�?                �]M�~a;�     �Y@                Y���@      "@     �7@��"��@        9����?�lscz�@�(�l*@        ����, �?�~j�t�J@:��7��@        �!XG���?      5@R��}
�@        ��ݮ��?                ��i�-(�      ;@                �7_w�z@      ,@n�2d�?#��Y%N@        @�H�{�?     �4@;�X��?        �E����?                Rl���+,@      .@                �bk++؞?      @]m�����?6�0�x @        ������?                        �k�g��?                85��@     @S@                vl�-�u@      4@                Qݾ
��      2@                w�1��      @                Qݾ
��      2@                w�1��      @     �>@�y)��E@              �?'�o|��?�	Ƹ�"@        �v���L�?5Sb�?3����M@        �D���Y�?��bb��?'�7�N@        ��]+'�?io����?99�%�*�?        XG��).�?                ʬ��c�5�     �S@                ׂ�b�!@     �S@                30�z��      S@                H�Q#3@     �L@                �^f�@      @                �J��@�@      @��� #@����@              �?8�9@��?�M��6@        Qj�a��?                        �k�g��?�H�}��?St�x��?        )5�0��?��Q���?�S2}*@        �Oq���?                �Ɵ� �1�     �[@                B��2@      g@:��K��?F4ש��@        J�=���?T���B�?��7���@        �}�K�`�?Z�����?                �k�g��?@x�=�?Lc�k@        �]+'<�?                �	�;ٞ3@     ``@                HZ~��#�     �J@Z�����?                XG��).�?���u�?�XO��A�?        �ߠ۵r�?                s?m��,@     @_@                HZ~��#�     �J@                ��>�@      3@                s�Φ7$@      c@                �Uws7�     �X@                �-\ӿ
@      @                ?d�W�
@      @                $@�y���      @      +@�qE@@              �?��E_A��?�̠�@	@        [9���?H�z�;@jwO�@        ���Y@��?                �)�a.�      G@                �&�t3�@      .@43333�6@f���|�@        )5�0ȧ?����̬E@����KQ�?        WNx��A�?                |'H��P@      "@                �.筟"@      @                ٮg��b�      A@                ��h�/ /@     �g@      /@'1_O�s@              �?      3@���!5
@        ��ݮ��?     @L@��i�@        �/���?                        ��ݮ��?     �<@QOk���?        �}�K�`�?                ���g0@     @m@                ������#�     �J@                ���g0@     @m@                ������#�     �J@                hUE�_@      @                hal+E	@      @      �?��2@              �?                        XG��).�?��� #@D�(@        �%C��6�?                ���\4�@      @                ���l��     pr@      #@w_����@        �/���?      B@[}I� @        �k�g��?�Բ�>�?j�"��?        @�H�{�?      @YN����@        Nx��A��?                q��JM�      @                ���C���      @                8酆�'�      9@                کv�i��?      @^�c@���?��pM�@        ��o��?      +@Xe�R@        �D���Y�?      <@A�p�\�@        &C��6�?     �?@e�V��@        �k�g��?3��V�?qW�A� @        ���:�?8�9@p�?����6@        t�VNx�?                ?瑖�.�     @[@                $�B����      @                �p�k~@     @S@                ��\jC)@      A@                �#x�R0@      4@                ��R��      @                �5��9�@      @                ,����	�      @1��*d�?-���(@              �?     �<@��2O@        .�u�y�?Z�8�ŭ�?                ;ڼOqɐ?      �?��4蹑@        1��R�?��Q��?@��UX�@        �t�VN�?                �nw0��4@     p@                �E <u�      B@                ����,m@      ,@                 ��;�%�     �e@                �؊/��@      @                ������0@      Y@      3@F�F��@              �?      @�*���} @        ާ�d��?     �8@�2QzY@        �����?                *�h��@      &@                7"��8�0�      Q@      '@��[���@        �k�g��?T��.q�?�lr�,@        ��E�Ը?                ���WG�      A@                yk�ƺ1@     �c@      C@�=e�&�?        �Y@�H��?      :@���D�?        j�a�/�?                r�I�@      @                 ��f@      @                ��)a��      @                I��J?@      0@��v��bO@��U~@              �?=
ףp�N@Uk��!�@        �, _$J�?�ʡE�#[@����D@        x��A�k�?                [�s�3�     �h@                X����      @                2�}�|(0@      W@                ��Y�L�      @��n��?��i�@              �?     �6@~�����@        ��|�(5�?��,`W@��~7�� @        ��ݮ��?      @��[8�T@        ��]+'�?      -@�du�"1@        h�t�V�?                �P�d'@      <@                ��W��@     �N@                        �"Qj�av?      -@,������?        �g�t�?�-�l�I�?>�ƅQ@        �D����?     �K@s.u�\@        v�y���?     �L@˽�^���?        �!XG��?*oG8-x�?                �/�Ǝ?      '@��ϮD @�"8��?      �?                        XG��).�?                ��^�4�4@      T@                ��0�d�      @                ٽ��R/�     �@@                ��$͟ �      ?@                �Zz�&�      G@                m�<?��?      @                Y$��d&�      H@                .�y��?      @                �H��#@       @                �f��d}&@      R@                �H��#@       @                �f��d}&@      R@      @�$J�^@              �?      �?_h��!��?        )5�0ȗ?     �D@^�yq8}@        WNx��A�?                �n�s��      @                �Lcǰ	�      @     �=@0��E�@        �u�y���?      +@��q�@        Sc��|�?                ��!bI *@     `d@                k#��|'�     �T@                ���ߟ�@      @                	�ɱ�"@     �C@      (@ыg%��@              �?                        �k�g�{?     �<@���� �@        )5�0��?                DEg�@      @                Ҩ��A�     �r@                UD]N`]2�      e@                z^��A�/@     �_@     �N@%^�W@              �?     @N@n�z���@        '<�ߠ��?     �a@�>j����?        �f�"�?     �8@���E��?        �, _$J�?                        j�a�/�?      #@�l�T�
@        @�H�{�?                        ��ݮ��?      @G�J �a@        Qj�a��?      J@�t����?        7�S\2�?                𹇱�J�?      b@                �-��J3@      `@X��0_��?_���*�?        )5�0ȗ?      '@ϖv��?        XG��).�?                �h��@      @                ]-y�,�?      &@                z �	U@      @                (�ەE�@      @                �*��      @                Ƶ|���?      @                �k[#]�@      @                ����.�     �a@                [�aZږ5@     �]@                �M�)�`�      "@     @J@�Q3�X@              �?     �R@⸖9GV@        �������?      '@��-�H�@        UUUUUU�?                Ҕ�1�@      l@                M}u�#@      6@                6��o]�0�     �C@                ɔ�Y$	@      (@     �G@yj
3@              �?��bٽ�?�9_�@        l�g��?     @J@�)�M�
@        )5�0��?     �R@�
�rv6@        8�v����?J$��(��?;�m/@        ?�%C���?                �u';�$�      3@                F�����     @U@     �]@��nP��@        ��o���?     0l@�\��l��?        #Qj�a�?                56�Lt�'�      =@                E���$�@      6@                ʝu� &@     �_@                Qx���@       @                9(�dG@      @                6��@      @                                �j�鳳?      �?      @      A@�"Qj�0@ �|!�w@               @      @     �Z@�, _$�@@���3@              @      @      P@ڼOq��7@ŵ+�)@              @        V�F�? @+�3X���?5��nݕ�?              @        ���4)@+���Č�?��v��]�?              @        rm���@z�����?��G�W�?              @        �zNz��@z�\�o�?���q?��?               @      "@     �d@}�(5��D@ub��C@              "@      "@      :@L�`m^0@v&��9�@              $@        \*���@����?sv���&�?              &@        Z����@>vVB+��?�G2���?              (@ףp=
W1@�(\��ug@����7R@�E�C@              *@        Nz���3
@t^Z:ZC�?��C$�v�?              ,@      $@     �r@2�h�NP@���%�O@              .@      9@      P@
��7��E@�p2�"@              0@      @      M@�g�t�;@��m�{\)@              1@      .@     �c@����I@���V7i:@              2@      @      =@F���ì-@�v�aH@              3@        ���V	V@[8<��O�?�$�j��?              4@       @     �M@��]+�5@�f�֗(@              5@        ��� E@����?��y����?              6@        ����%@=�^���?{|��5[�?              7@        H�I�O��?`a�x���?�Ì,���?              8@       @      .@
��7�v@��c�/@              9@      @      3@�H�{�!@P�z�a@              :@      @      6@�:ڼO�$@��/.�O@              ;@       @      V@*.�uA@_��c�1@              <@      @      .@�o��Z9!@U�v�@              =@        [닄�\@I����?�.H��h�?              >@        AJ�i;	@iu�#��?�#u!h�?              ?@             �M@���.9@����-@              @@       @      9@��6�S\&@*J��X�@             �@@       @      @@�y��!3@��11��@              A@        ;�f�_ @�~��uK�?���>�� @             �A@        �D�
)� @N;J��*�?�tL�s @              B@      1@     0u@��}�K&P@]y��(�M@             �B@      �?      ?@��f�*@�r*h��@              C@        �����@e/ٻ�\�?]v��0��?             �C@              b@�7�v��J@�W)�B@              D@              M@4��]+5@K��� �*@             �D@        �SW>+@�(�|E�?\�����?              E@{�G��3@ףp=
\@f�k��3L@�,I�xi6@             �E@        ��.�@g��k�?�a�����?              F@      *@     �r@�r�3�I@��>Ai$J@             �F@        |a2U0�?CB�����?舎e�?              G@        ���K�@�Bq�t�?v%'���?             �G@        %̴�+�@z0��L�?��D���?              H@        �@+0du�?itq	S��?sJ� 6�?             �H@       @      ;@�}�K�`0@�`P�@              I@        �����@E/]t��?�S|�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        